// File:    jpeg_tb.sv
// Author:  Lei Kuang
// Date:    17th June 2020
// @ Imperial College London

module jpeg_tb;

logic        clk;
logic        nrst;
logic [7:0]  din;
logic        din_valid;
logic [31:0] dout;
logic        dout_valid;

jpeg dut(.*);

initial begin
    clk = '0;
    forever #5ns clk = ~clk;
end

logic [13:0] din_cnt;
logic [7:0]  img [16383:0];

logic [7:0] cnt;

initial begin
    cnt = '0;
    
    @(posedge nrst)
    ;
    
    forever @ (posedge clk)
        cnt = cnt + 1;
end

assign din_valid = cnt=='1;

initial begin
    nrst      = '0;
    din_cnt   = '0;
    
    @(posedge clk)
        nrst <= '1;
    
    forever begin
        @(posedge clk) begin
            if(din_valid)
                din_cnt <= din_cnt + 1;
        end
    end
end

assign din = img[din_cnt];

initial begin
    forever @ (negedge clk) begin
        if(dout_valid)
            $write("%X\n", dout);
    end
end

// img = plt.imread('./blackpearl/bmp/batman_1.bmp', 0)
begin
assign img[    0] = 0;
assign img[    1] = 204;
assign img[    2] = 236;
assign img[    3] = 238;
assign img[    4] = 238;
assign img[    5] = 238;
assign img[    6] = 206;
assign img[    7] = 238;
assign img[    8] = 254;
assign img[    9] = 255;
assign img[   10] = 255;
assign img[   11] = 239;
assign img[   12] = 204;
assign img[   13] = 236;
assign img[   14] = 238;
assign img[   15] = 191;
assign img[   16] = 187;
assign img[   17] = 239;
assign img[   18] = 238;
assign img[   19] = 174;
assign img[   20] = 170;
assign img[   21] = 238;
assign img[   22] = 238;
assign img[   23] = 238;
assign img[   24] = 238;
assign img[   25] = 238;
assign img[   26] = 204;
assign img[   27] = 236;
assign img[   28] = 206;
assign img[   29] = 236;
assign img[   30] = 238;
assign img[   31] = 255;
assign img[   32] = 239;
assign img[   33] = 238;
assign img[   34] = 254;
assign img[   35] = 255;
assign img[   36] = 255;
assign img[   37] = 255;
assign img[   38] = 254;
assign img[   39] = 255;
assign img[   40] = 238;
assign img[   41] = 238;
assign img[   42] = 238;
assign img[   43] = 238;
assign img[   44] = 238;
assign img[   45] = 254;
assign img[   46] = 255;
assign img[   47] = 255;
assign img[   48] = 255;
assign img[   49] = 255;
assign img[   50] = 223;
assign img[   51] = 255;
assign img[   52] = 255;
assign img[   53] = 255;
assign img[   54] = 255;
assign img[   55] = 255;
assign img[   56] = 255;
assign img[   57] = 255;
assign img[   58] = 255;
assign img[   59] = 255;
assign img[   60] = 238;
assign img[   61] = 238;
assign img[   62] = 238;
assign img[   63] = 255;
assign img[   64] = 255;
assign img[   65] = 255;
assign img[   66] = 255;
assign img[   67] = 255;
assign img[   68] = 255;
assign img[   69] = 255;
assign img[   70] = 221;
assign img[   71] = 239;
assign img[   72] = 238;
assign img[   73] = 238;
assign img[   74] = 254;
assign img[   75] = 239;
assign img[   76] = 238;
assign img[   77] = 223;
assign img[   78] = 255;
assign img[   79] = 255;
assign img[   80] = 223;
assign img[   81] = 255;
assign img[   82] = 255;
assign img[   83] = 255;
assign img[   84] = 238;
assign img[   85] = 255;
assign img[   86] = 255;
assign img[   87] = 255;
assign img[   88] = 239;
assign img[   89] = 255;
assign img[   90] = 255;
assign img[   91] = 255;
assign img[   92] = 255;
assign img[   93] = 255;
assign img[   94] = 254;
assign img[   95] = 191;
assign img[   96] = 170;
assign img[   97] = 234;
assign img[   98] = 238;
assign img[   99] = 142;
assign img[  100] = 238;
assign img[  101] = 255;
assign img[  102] = 221;
assign img[  103] = 253;
assign img[  104] = 238;
assign img[  105] = 255;
assign img[  106] = 255;
assign img[  107] = 239;
assign img[  108] = 206;
assign img[  109] = 238;
assign img[  110] = 238;
assign img[  111] = 254;
assign img[  112] = 221;
assign img[  113] = 255;
assign img[  114] = 255;
assign img[  115] = 255;
assign img[  116] = 221;
assign img[  117] = 253;
assign img[  118] = 255;
assign img[  119] = 223;
assign img[  120] = 221;
assign img[  121] = 221;
assign img[  122] = 253;
assign img[  123] = 255;
assign img[  124] = 255;
assign img[  125] = 255;
assign img[  126] = 255;
assign img[  127] = 255;
assign img[  128] = 96;
assign img[  129] = 238;
assign img[  130] = 238;
assign img[  131] = 255;
assign img[  132] = 255;
assign img[  133] = 255;
assign img[  134] = 191;
assign img[  135] = 238;
assign img[  136] = 238;
assign img[  137] = 255;
assign img[  138] = 254;
assign img[  139] = 238;
assign img[  140] = 238;
assign img[  141] = 238;
assign img[  142] = 238;
assign img[  143] = 238;
assign img[  144] = 204;
assign img[  145] = 204;
assign img[  146] = 238;
assign img[  147] = 255;
assign img[  148] = 238;
assign img[  149] = 255;
assign img[  150] = 255;
assign img[  151] = 255;
assign img[  152] = 255;
assign img[  153] = 255;
assign img[  154] = 138;
assign img[  155] = 238;
assign img[  156] = 238;
assign img[  157] = 255;
assign img[  158] = 239;
assign img[  159] = 206;
assign img[  160] = 236;
assign img[  161] = 238;
assign img[  162] = 238;
assign img[  163] = 238;
assign img[  164] = 238;
assign img[  165] = 238;
assign img[  166] = 254;
assign img[  167] = 223;
assign img[  168] = 253;
assign img[  169] = 255;
assign img[  170] = 239;
assign img[  171] = 238;
assign img[  172] = 238;
assign img[  173] = 239;
assign img[  174] = 238;
assign img[  175] = 255;
assign img[  176] = 255;
assign img[  177] = 255;
assign img[  178] = 255;
assign img[  179] = 255;
assign img[  180] = 255;
assign img[  181] = 255;
assign img[  182] = 255;
assign img[  183] = 255;
assign img[  184] = 255;
assign img[  185] = 255;
assign img[  186] = 239;
assign img[  187] = 254;
assign img[  188] = 255;
assign img[  189] = 255;
assign img[  190] = 255;
assign img[  191] = 255;
assign img[  192] = 255;
assign img[  193] = 255;
assign img[  194] = 255;
assign img[  195] = 255;
assign img[  196] = 255;
assign img[  197] = 255;
assign img[  198] = 238;
assign img[  199] = 238;
assign img[  200] = 238;
assign img[  201] = 255;
assign img[  202] = 255;
assign img[  203] = 223;
assign img[  204] = 255;
assign img[  205] = 255;
assign img[  206] = 255;
assign img[  207] = 255;
assign img[  208] = 255;
assign img[  209] = 255;
assign img[  210] = 239;
assign img[  211] = 238;
assign img[  212] = 238;
assign img[  213] = 207;
assign img[  214] = 236;
assign img[  215] = 238;
assign img[  216] = 238;
assign img[  217] = 255;
assign img[  218] = 223;
assign img[  219] = 221;
assign img[  220] = 236;
assign img[  221] = 238;
assign img[  222] = 238;
assign img[  223] = 174;
assign img[  224] = 238;
assign img[  225] = 238;
assign img[  226] = 254;
assign img[  227] = 255;
assign img[  228] = 255;
assign img[  229] = 207;
assign img[  230] = 204;
assign img[  231] = 254;
assign img[  232] = 255;
assign img[  233] = 255;
assign img[  234] = 238;
assign img[  235] = 238;
assign img[  236] = 206;
assign img[  237] = 238;
assign img[  238] = 238;
assign img[  239] = 238;
assign img[  240] = 238;
assign img[  241] = 238;
assign img[  242] = 238;
assign img[  243] = 238;
assign img[  244] = 254;
assign img[  245] = 255;
assign img[  246] = 238;
assign img[  247] = 239;
assign img[  248] = 254;
assign img[  249] = 238;
assign img[  250] = 238;
assign img[  251] = 255;
assign img[  252] = 221;
assign img[  253] = 253;
assign img[  254] = 255;
assign img[  255] = 255;
assign img[  256] = 96;
assign img[  257] = 238;
assign img[  258] = 238;
assign img[  259] = 238;
assign img[  260] = 186;
assign img[  261] = 251;
assign img[  262] = 239;
assign img[  263] = 254;
assign img[  264] = 255;
assign img[  265] = 255;
assign img[  266] = 255;
assign img[  267] = 255;
assign img[  268] = 221;
assign img[  269] = 255;
assign img[  270] = 255;
assign img[  271] = 255;
assign img[  272] = 204;
assign img[  273] = 254;
assign img[  274] = 254;
assign img[  275] = 238;
assign img[  276] = 254;
assign img[  277] = 255;
assign img[  278] = 255;
assign img[  279] = 255;
assign img[  280] = 238;
assign img[  281] = 255;
assign img[  282] = 255;
assign img[  283] = 255;
assign img[  284] = 255;
assign img[  285] = 255;
assign img[  286] = 255;
assign img[  287] = 191;
assign img[  288] = 255;
assign img[  289] = 255;
assign img[  290] = 255;
assign img[  291] = 255;
assign img[  292] = 255;
assign img[  293] = 255;
assign img[  294] = 255;
assign img[  295] = 255;
assign img[  296] = 255;
assign img[  297] = 255;
assign img[  298] = 255;
assign img[  299] = 239;
assign img[  300] = 238;
assign img[  301] = 238;
assign img[  302] = 238;
assign img[  303] = 255;
assign img[  304] = 255;
assign img[  305] = 255;
assign img[  306] = 255;
assign img[  307] = 255;
assign img[  308] = 255;
assign img[  309] = 255;
assign img[  310] = 255;
assign img[  311] = 255;
assign img[  312] = 255;
assign img[  313] = 239;
assign img[  314] = 222;
assign img[  315] = 221;
assign img[  316] = 253;
assign img[  317] = 255;
assign img[  318] = 223;
assign img[  319] = 253;
assign img[  320] = 255;
assign img[  321] = 223;
assign img[  322] = 238;
assign img[  323] = 238;
assign img[  324] = 222;
assign img[  325] = 223;
assign img[  326] = 255;
assign img[  327] = 238;
assign img[  328] = 238;
assign img[  329] = 238;
assign img[  330] = 255;
assign img[  331] = 255;
assign img[  332] = 255;
assign img[  333] = 255;
assign img[  334] = 255;
assign img[  335] = 255;
assign img[  336] = 255;
assign img[  337] = 255;
assign img[  338] = 255;
assign img[  339] = 255;
assign img[  340] = 223;
assign img[  341] = 221;
assign img[  342] = 253;
assign img[  343] = 255;
assign img[  344] = 255;
assign img[  345] = 255;
assign img[  346] = 255;
assign img[  347] = 239;
assign img[  348] = 238;
assign img[  349] = 238;
assign img[  350] = 238;
assign img[  351] = 255;
assign img[  352] = 255;
assign img[  353] = 255;
assign img[  354] = 255;
assign img[  355] = 255;
assign img[  356] = 255;
assign img[  357] = 239;
assign img[  358] = 238;
assign img[  359] = 238;
assign img[  360] = 238;
assign img[  361] = 255;
assign img[  362] = 255;
assign img[  363] = 255;
assign img[  364] = 255;
assign img[  365] = 255;
assign img[  366] = 255;
assign img[  367] = 255;
assign img[  368] = 255;
assign img[  369] = 255;
assign img[  370] = 255;
assign img[  371] = 239;
assign img[  372] = 238;
assign img[  373] = 238;
assign img[  374] = 238;
assign img[  375] = 238;
assign img[  376] = 238;
assign img[  377] = 255;
assign img[  378] = 238;
assign img[  379] = 174;
assign img[  380] = 186;
assign img[  381] = 251;
assign img[  382] = 255;
assign img[  383] = 255;
assign img[  384] = 96;
assign img[  385] = 238;
assign img[  386] = 238;
assign img[  387] = 239;
assign img[  388] = 238;
assign img[  389] = 238;
assign img[  390] = 254;
assign img[  391] = 223;
assign img[  392] = 253;
assign img[  393] = 255;
assign img[  394] = 255;
assign img[  395] = 255;
assign img[  396] = 221;
assign img[  397] = 253;
assign img[  398] = 255;
assign img[  399] = 223;
assign img[  400] = 204;
assign img[  401] = 204;
assign img[  402] = 238;
assign img[  403] = 239;
assign img[  404] = 186;
assign img[  405] = 238;
assign img[  406] = 255;
assign img[  407] = 255;
assign img[  408] = 255;
assign img[  409] = 191;
assign img[  410] = 187;
assign img[  411] = 255;
assign img[  412] = 255;
assign img[  413] = 255;
assign img[  414] = 255;
assign img[  415] = 239;
assign img[  416] = 78;
assign img[  417] = 255;
assign img[  418] = 255;
assign img[  419] = 255;
assign img[  420] = 191;
assign img[  421] = 187;
assign img[  422] = 251;
assign img[  423] = 255;
assign img[  424] = 255;
assign img[  425] = 255;
assign img[  426] = 239;
assign img[  427] = 238;
assign img[  428] = 238;
assign img[  429] = 239;
assign img[  430] = 238;
assign img[  431] = 238;
assign img[  432] = 254;
assign img[  433] = 255;
assign img[  434] = 255;
assign img[  435] = 255;
assign img[  436] = 238;
assign img[  437] = 238;
assign img[  438] = 222;
assign img[  439] = 255;
assign img[  440] = 255;
assign img[  441] = 223;
assign img[  442] = 205;
assign img[  443] = 238;
assign img[  444] = 238;
assign img[  445] = 175;
assign img[  446] = 238;
assign img[  447] = 238;
assign img[  448] = 238;
assign img[  449] = 238;
assign img[  450] = 174;
assign img[  451] = 238;
assign img[  452] = 238;
assign img[  453] = 254;
assign img[  454] = 255;
assign img[  455] = 255;
assign img[  456] = 238;
assign img[  457] = 255;
assign img[  458] = 255;
assign img[  459] = 255;
assign img[  460] = 239;
assign img[  461] = 238;
assign img[  462] = 238;
assign img[  463] = 255;
assign img[  464] = 255;
assign img[  465] = 255;
assign img[  466] = 255;
assign img[  467] = 255;
assign img[  468] = 255;
assign img[  469] = 255;
assign img[  470] = 238;
assign img[  471] = 238;
assign img[  472] = 238;
assign img[  473] = 238;
assign img[  474] = 238;
assign img[  475] = 191;
assign img[  476] = 251;
assign img[  477] = 255;
assign img[  478] = 255;
assign img[  479] = 223;
assign img[  480] = 221;
assign img[  481] = 205;
assign img[  482] = 252;
assign img[  483] = 255;
assign img[  484] = 255;
assign img[  485] = 239;
assign img[  486] = 204;
assign img[  487] = 238;
assign img[  488] = 238;
assign img[  489] = 238;
assign img[  490] = 238;
assign img[  491] = 255;
assign img[  492] = 238;
assign img[  493] = 238;
assign img[  494] = 238;
assign img[  495] = 254;
assign img[  496] = 223;
assign img[  497] = 221;
assign img[  498] = 253;
assign img[  499] = 255;
assign img[  500] = 204;
assign img[  501] = 253;
assign img[  502] = 255;
assign img[  503] = 255;
assign img[  504] = 223;
assign img[  505] = 255;
assign img[  506] = 187;
assign img[  507] = 223;
assign img[  508] = 221;
assign img[  509] = 255;
assign img[  510] = 255;
assign img[  511] = 255;
assign img[  512] = 96;
assign img[  513] = 238;
assign img[  514] = 254;
assign img[  515] = 255;
assign img[  516] = 223;
assign img[  517] = 221;
assign img[  518] = 253;
assign img[  519] = 254;
assign img[  520] = 238;
assign img[  521] = 255;
assign img[  522] = 254;
assign img[  523] = 238;
assign img[  524] = 220;
assign img[  525] = 253;
assign img[  526] = 255;
assign img[  527] = 255;
assign img[  528] = 221;
assign img[  529] = 253;
assign img[  530] = 255;
assign img[  531] = 223;
assign img[  532] = 221;
assign img[  533] = 253;
assign img[  534] = 255;
assign img[  535] = 255;
assign img[  536] = 255;
assign img[  537] = 239;
assign img[  538] = 238;
assign img[  539] = 238;
assign img[  540] = 238;
assign img[  541] = 238;
assign img[  542] = 254;
assign img[  543] = 207;
assign img[  544] = 204;
assign img[  545] = 238;
assign img[  546] = 238;
assign img[  547] = 238;
assign img[  548] = 238;
assign img[  549] = 239;
assign img[  550] = 206;
assign img[  551] = 204;
assign img[  552] = 236;
assign img[  553] = 238;
assign img[  554] = 206;
assign img[  555] = 238;
assign img[  556] = 222;
assign img[  557] = 221;
assign img[  558] = 253;
assign img[  559] = 239;
assign img[  560] = 254;
assign img[  561] = 255;
assign img[  562] = 255;
assign img[  563] = 255;
assign img[  564] = 255;
assign img[  565] = 255;
assign img[  566] = 255;
assign img[  567] = 255;
assign img[  568] = 255;
assign img[  569] = 255;
assign img[  570] = 255;
assign img[  571] = 255;
assign img[  572] = 255;
assign img[  573] = 255;
assign img[  574] = 221;
assign img[  575] = 253;
assign img[  576] = 255;
assign img[  577] = 223;
assign img[  578] = 205;
assign img[  579] = 236;
assign img[  580] = 254;
assign img[  581] = 255;
assign img[  582] = 255;
assign img[  583] = 255;
assign img[  584] = 255;
assign img[  585] = 239;
assign img[  586] = 254;
assign img[  587] = 255;
assign img[  588] = 239;
assign img[  589] = 238;
assign img[  590] = 238;
assign img[  591] = 255;
assign img[  592] = 255;
assign img[  593] = 255;
assign img[  594] = 255;
assign img[  595] = 223;
assign img[  596] = 253;
assign img[  597] = 255;
assign img[  598] = 238;
assign img[  599] = 238;
assign img[  600] = 206;
assign img[  601] = 220;
assign img[  602] = 237;
assign img[  603] = 238;
assign img[  604] = 238;
assign img[  605] = 238;
assign img[  606] = 238;
assign img[  607] = 206;
assign img[  608] = 238;
assign img[  609] = 204;
assign img[  610] = 238;
assign img[  611] = 238;
assign img[  612] = 238;
assign img[  613] = 255;
assign img[  614] = 221;
assign img[  615] = 255;
assign img[  616] = 238;
assign img[  617] = 254;
assign img[  618] = 238;
assign img[  619] = 255;
assign img[  620] = 221;
assign img[  621] = 253;
assign img[  622] = 255;
assign img[  623] = 223;
assign img[  624] = 221;
assign img[  625] = 253;
assign img[  626] = 255;
assign img[  627] = 255;
assign img[  628] = 221;
assign img[  629] = 253;
assign img[  630] = 255;
assign img[  631] = 255;
assign img[  632] = 255;
assign img[  633] = 239;
assign img[  634] = 238;
assign img[  635] = 254;
assign img[  636] = 255;
assign img[  637] = 255;
assign img[  638] = 255;
assign img[  639] = 255;
assign img[  640] = 96;
assign img[  641] = 238;
assign img[  642] = 238;
assign img[  643] = 206;
assign img[  644] = 204;
assign img[  645] = 252;
assign img[  646] = 206;
assign img[  647] = 236;
assign img[  648] = 238;
assign img[  649] = 238;
assign img[  650] = 254;
assign img[  651] = 239;
assign img[  652] = 238;
assign img[  653] = 254;
assign img[  654] = 255;
assign img[  655] = 191;
assign img[  656] = 187;
assign img[  657] = 251;
assign img[  658] = 238;
assign img[  659] = 255;
assign img[  660] = 255;
assign img[  661] = 255;
assign img[  662] = 238;
assign img[  663] = 254;
assign img[  664] = 239;
assign img[  665] = 238;
assign img[  666] = 238;
assign img[  667] = 238;
assign img[  668] = 238;
assign img[  669] = 238;
assign img[  670] = 238;
assign img[  671] = 174;
assign img[  672] = 220;
assign img[  673] = 255;
assign img[  674] = 255;
assign img[  675] = 255;
assign img[  676] = 255;
assign img[  677] = 255;
assign img[  678] = 255;
assign img[  679] = 255;
assign img[  680] = 255;
assign img[  681] = 255;
assign img[  682] = 255;
assign img[  683] = 255;
assign img[  684] = 255;
assign img[  685] = 255;
assign img[  686] = 238;
assign img[  687] = 255;
assign img[  688] = 255;
assign img[  689] = 255;
assign img[  690] = 255;
assign img[  691] = 255;
assign img[  692] = 255;
assign img[  693] = 255;
assign img[  694] = 255;
assign img[  695] = 255;
assign img[  696] = 255;
assign img[  697] = 255;
assign img[  698] = 255;
assign img[  699] = 255;
assign img[  700] = 255;
assign img[  701] = 238;
assign img[  702] = 238;
assign img[  703] = 255;
assign img[  704] = 255;
assign img[  705] = 255;
assign img[  706] = 255;
assign img[  707] = 255;
assign img[  708] = 255;
assign img[  709] = 239;
assign img[  710] = 238;
assign img[  711] = 238;
assign img[  712] = 238;
assign img[  713] = 238;
assign img[  714] = 238;
assign img[  715] = 254;
assign img[  716] = 238;
assign img[  717] = 238;
assign img[  718] = 238;
assign img[  719] = 255;
assign img[  720] = 223;
assign img[  721] = 255;
assign img[  722] = 239;
assign img[  723] = 238;
assign img[  724] = 238;
assign img[  725] = 238;
assign img[  726] = 238;
assign img[  727] = 238;
assign img[  728] = 206;
assign img[  729] = 254;
assign img[  730] = 255;
assign img[  731] = 255;
assign img[  732] = 255;
assign img[  733] = 255;
assign img[  734] = 255;
assign img[  735] = 255;
assign img[  736] = 187;
assign img[  737] = 251;
assign img[  738] = 255;
assign img[  739] = 255;
assign img[  740] = 255;
assign img[  741] = 255;
assign img[  742] = 191;
assign img[  743] = 255;
assign img[  744] = 255;
assign img[  745] = 255;
assign img[  746] = 238;
assign img[  747] = 254;
assign img[  748] = 175;
assign img[  749] = 255;
assign img[  750] = 238;
assign img[  751] = 174;
assign img[  752] = 170;
assign img[  753] = 170;
assign img[  754] = 234;
assign img[  755] = 238;
assign img[  756] = 239;
assign img[  757] = 255;
assign img[  758] = 255;
assign img[  759] = 255;
assign img[  760] = 255;
assign img[  761] = 255;
assign img[  762] = 238;
assign img[  763] = 238;
assign img[  764] = 220;
assign img[  765] = 253;
assign img[  766] = 255;
assign img[  767] = 255;
assign img[  768] = 96;
assign img[  769] = 238;
assign img[  770] = 254;
assign img[  771] = 255;
assign img[  772] = 238;
assign img[  773] = 238;
assign img[  774] = 254;
assign img[  775] = 255;
assign img[  776] = 255;
assign img[  777] = 255;
assign img[  778] = 254;
assign img[  779] = 223;
assign img[  780] = 253;
assign img[  781] = 255;
assign img[  782] = 223;
assign img[  783] = 221;
assign img[  784] = 253;
assign img[  785] = 255;
assign img[  786] = 255;
assign img[  787] = 191;
assign img[  788] = 187;
assign img[  789] = 255;
assign img[  790] = 255;
assign img[  791] = 255;
assign img[  792] = 255;
assign img[  793] = 255;
assign img[  794] = 221;
assign img[  795] = 255;
assign img[  796] = 255;
assign img[  797] = 255;
assign img[  798] = 255;
assign img[  799] = 255;
assign img[  800] = 238;
assign img[  801] = 238;
assign img[  802] = 238;
assign img[  803] = 238;
assign img[  804] = 254;
assign img[  805] = 255;
assign img[  806] = 255;
assign img[  807] = 255;
assign img[  808] = 255;
assign img[  809] = 255;
assign img[  810] = 223;
assign img[  811] = 239;
assign img[  812] = 238;
assign img[  813] = 255;
assign img[  814] = 255;
assign img[  815] = 255;
assign img[  816] = 255;
assign img[  817] = 255;
assign img[  818] = 255;
assign img[  819] = 239;
assign img[  820] = 238;
assign img[  821] = 238;
assign img[  822] = 238;
assign img[  823] = 238;
assign img[  824] = 238;
assign img[  825] = 238;
assign img[  826] = 238;
assign img[  827] = 254;
assign img[  828] = 255;
assign img[  829] = 255;
assign img[  830] = 239;
assign img[  831] = 255;
assign img[  832] = 255;
assign img[  833] = 223;
assign img[  834] = 204;
assign img[  835] = 236;
assign img[  836] = 255;
assign img[  837] = 239;
assign img[  838] = 238;
assign img[  839] = 238;
assign img[  840] = 254;
assign img[  841] = 255;
assign img[  842] = 255;
assign img[  843] = 239;
assign img[  844] = 238;
assign img[  845] = 238;
assign img[  846] = 238;
assign img[  847] = 255;
assign img[  848] = 223;
assign img[  849] = 255;
assign img[  850] = 255;
assign img[  851] = 255;
assign img[  852] = 255;
assign img[  853] = 255;
assign img[  854] = 255;
assign img[  855] = 255;
assign img[  856] = 255;
assign img[  857] = 255;
assign img[  858] = 255;
assign img[  859] = 255;
assign img[  860] = 255;
assign img[  861] = 255;
assign img[  862] = 255;
assign img[  863] = 191;
assign img[  864] = 138;
assign img[  865] = 238;
assign img[  866] = 254;
assign img[  867] = 255;
assign img[  868] = 255;
assign img[  869] = 239;
assign img[  870] = 238;
assign img[  871] = 238;
assign img[  872] = 238;
assign img[  873] = 255;
assign img[  874] = 255;
assign img[  875] = 255;
assign img[  876] = 255;
assign img[  877] = 255;
assign img[  878] = 255;
assign img[  879] = 255;
assign img[  880] = 255;
assign img[  881] = 255;
assign img[  882] = 255;
assign img[  883] = 239;
assign img[  884] = 222;
assign img[  885] = 255;
assign img[  886] = 255;
assign img[  887] = 255;
assign img[  888] = 255;
assign img[  889] = 255;
assign img[  890] = 255;
assign img[  891] = 255;
assign img[  892] = 238;
assign img[  893] = 254;
assign img[  894] = 255;
assign img[  895] = 255;
assign img[  896] = 0;
assign img[  897] = 204;
assign img[  898] = 236;
assign img[  899] = 238;
assign img[  900] = 204;
assign img[  901] = 204;
assign img[  902] = 204;
assign img[  903] = 204;
assign img[  904] = 236;
assign img[  905] = 238;
assign img[  906] = 238;
assign img[  907] = 223;
assign img[  908] = 205;
assign img[  909] = 236;
assign img[  910] = 222;
assign img[  911] = 205;
assign img[  912] = 220;
assign img[  913] = 221;
assign img[  914] = 255;
assign img[  915] = 191;
assign img[  916] = 187;
assign img[  917] = 255;
assign img[  918] = 191;
assign img[  919] = 255;
assign img[  920] = 255;
assign img[  921] = 239;
assign img[  922] = 204;
assign img[  923] = 236;
assign img[  924] = 238;
assign img[  925] = 255;
assign img[  926] = 255;
assign img[  927] = 255;
assign img[  928] = 238;
assign img[  929] = 255;
assign img[  930] = 255;
assign img[  931] = 255;
assign img[  932] = 255;
assign img[  933] = 239;
assign img[  934] = 254;
assign img[  935] = 255;
assign img[  936] = 205;
assign img[  937] = 236;
assign img[  938] = 238;
assign img[  939] = 238;
assign img[  940] = 238;
assign img[  941] = 239;
assign img[  942] = 238;
assign img[  943] = 255;
assign img[  944] = 255;
assign img[  945] = 255;
assign img[  946] = 255;
assign img[  947] = 239;
assign img[  948] = 238;
assign img[  949] = 255;
assign img[  950] = 255;
assign img[  951] = 255;
assign img[  952] = 255;
assign img[  953] = 255;
assign img[  954] = 223;
assign img[  955] = 255;
assign img[  956] = 255;
assign img[  957] = 255;
assign img[  958] = 238;
assign img[  959] = 255;
assign img[  960] = 255;
assign img[  961] = 255;
assign img[  962] = 239;
assign img[  963] = 238;
assign img[  964] = 238;
assign img[  965] = 238;
assign img[  966] = 238;
assign img[  967] = 238;
assign img[  968] = 238;
assign img[  969] = 238;
assign img[  970] = 254;
assign img[  971] = 255;
assign img[  972] = 255;
assign img[  973] = 255;
assign img[  974] = 255;
assign img[  975] = 255;
assign img[  976] = 239;
assign img[  977] = 238;
assign img[  978] = 238;
assign img[  979] = 238;
assign img[  980] = 238;
assign img[  981] = 238;
assign img[  982] = 238;
assign img[  983] = 239;
assign img[  984] = 238;
assign img[  985] = 255;
assign img[  986] = 255;
assign img[  987] = 255;
assign img[  988] = 255;
assign img[  989] = 255;
assign img[  990] = 255;
assign img[  991] = 191;
assign img[  992] = 171;
assign img[  993] = 238;
assign img[  994] = 254;
assign img[  995] = 255;
assign img[  996] = 255;
assign img[  997] = 255;
assign img[  998] = 221;
assign img[  999] = 253;
assign img[ 1000] = 255;
assign img[ 1001] = 255;
assign img[ 1002] = 255;
assign img[ 1003] = 255;
assign img[ 1004] = 255;
assign img[ 1005] = 255;
assign img[ 1006] = 239;
assign img[ 1007] = 206;
assign img[ 1008] = 204;
assign img[ 1009] = 206;
assign img[ 1010] = 254;
assign img[ 1011] = 207;
assign img[ 1012] = 204;
assign img[ 1013] = 221;
assign img[ 1014] = 253;
assign img[ 1015] = 255;
assign img[ 1016] = 255;
assign img[ 1017] = 255;
assign img[ 1018] = 238;
assign img[ 1019] = 238;
assign img[ 1020] = 238;
assign img[ 1021] = 238;
assign img[ 1022] = 254;
assign img[ 1023] = 223;
assign img[ 1024] = 96;
assign img[ 1025] = 239;
assign img[ 1026] = 238;
assign img[ 1027] = 223;
assign img[ 1028] = 205;
assign img[ 1029] = 252;
assign img[ 1030] = 221;
assign img[ 1031] = 221;
assign img[ 1032] = 236;
assign img[ 1033] = 223;
assign img[ 1034] = 157;
assign img[ 1035] = 136;
assign img[ 1036] = 200;
assign img[ 1037] = 204;
assign img[ 1038] = 220;
assign img[ 1039] = 221;
assign img[ 1040] = 255;
assign img[ 1041] = 255;
assign img[ 1042] = 254;
assign img[ 1043] = 255;
assign img[ 1044] = 239;
assign img[ 1045] = 238;
assign img[ 1046] = 238;
assign img[ 1047] = 238;
assign img[ 1048] = 238;
assign img[ 1049] = 255;
assign img[ 1050] = 187;
assign img[ 1051] = 251;
assign img[ 1052] = 255;
assign img[ 1053] = 255;
assign img[ 1054] = 239;
assign img[ 1055] = 206;
assign img[ 1056] = 236;
assign img[ 1057] = 255;
assign img[ 1058] = 175;
assign img[ 1059] = 254;
assign img[ 1060] = 239;
assign img[ 1061] = 238;
assign img[ 1062] = 254;
assign img[ 1063] = 255;
assign img[ 1064] = 255;
assign img[ 1065] = 255;
assign img[ 1066] = 255;
assign img[ 1067] = 255;
assign img[ 1068] = 238;
assign img[ 1069] = 238;
assign img[ 1070] = 238;
assign img[ 1071] = 255;
assign img[ 1072] = 238;
assign img[ 1073] = 238;
assign img[ 1074] = 238;
assign img[ 1075] = 255;
assign img[ 1076] = 255;
assign img[ 1077] = 255;
assign img[ 1078] = 255;
assign img[ 1079] = 255;
assign img[ 1080] = 223;
assign img[ 1081] = 221;
assign img[ 1082] = 221;
assign img[ 1083] = 255;
assign img[ 1084] = 255;
assign img[ 1085] = 255;
assign img[ 1086] = 255;
assign img[ 1087] = 255;
assign img[ 1088] = 255;
assign img[ 1089] = 255;
assign img[ 1090] = 239;
assign img[ 1091] = 255;
assign img[ 1092] = 255;
assign img[ 1093] = 239;
assign img[ 1094] = 238;
assign img[ 1095] = 238;
assign img[ 1096] = 238;
assign img[ 1097] = 255;
assign img[ 1098] = 255;
assign img[ 1099] = 255;
assign img[ 1100] = 255;
assign img[ 1101] = 255;
assign img[ 1102] = 255;
assign img[ 1103] = 255;
assign img[ 1104] = 239;
assign img[ 1105] = 238;
assign img[ 1106] = 222;
assign img[ 1107] = 255;
assign img[ 1108] = 239;
assign img[ 1109] = 238;
assign img[ 1110] = 238;
assign img[ 1111] = 238;
assign img[ 1112] = 238;
assign img[ 1113] = 255;
assign img[ 1114] = 255;
assign img[ 1115] = 255;
assign img[ 1116] = 255;
assign img[ 1117] = 255;
assign img[ 1118] = 255;
assign img[ 1119] = 191;
assign img[ 1120] = 251;
assign img[ 1121] = 255;
assign img[ 1122] = 255;
assign img[ 1123] = 255;
assign img[ 1124] = 255;
assign img[ 1125] = 223;
assign img[ 1126] = 237;
assign img[ 1127] = 238;
assign img[ 1128] = 238;
assign img[ 1129] = 238;
assign img[ 1130] = 238;
assign img[ 1131] = 239;
assign img[ 1132] = 238;
assign img[ 1133] = 238;
assign img[ 1134] = 238;
assign img[ 1135] = 238;
assign img[ 1136] = 255;
assign img[ 1137] = 255;
assign img[ 1138] = 239;
assign img[ 1139] = 206;
assign img[ 1140] = 204;
assign img[ 1141] = 174;
assign img[ 1142] = 138;
assign img[ 1143] = 236;
assign img[ 1144] = 238;
assign img[ 1145] = 238;
assign img[ 1146] = 204;
assign img[ 1147] = 204;
assign img[ 1148] = 204;
assign img[ 1149] = 236;
assign img[ 1150] = 238;
assign img[ 1151] = 238;
assign img[ 1152] = 96;
assign img[ 1153] = 159;
assign img[ 1154] = 249;
assign img[ 1155] = 255;
assign img[ 1156] = 221;
assign img[ 1157] = 221;
assign img[ 1158] = 253;
assign img[ 1159] = 255;
assign img[ 1160] = 255;
assign img[ 1161] = 255;
assign img[ 1162] = 255;
assign img[ 1163] = 255;
assign img[ 1164] = 255;
assign img[ 1165] = 255;
assign img[ 1166] = 239;
assign img[ 1167] = 238;
assign img[ 1168] = 238;
assign img[ 1169] = 238;
assign img[ 1170] = 238;
assign img[ 1171] = 174;
assign img[ 1172] = 170;
assign img[ 1173] = 238;
assign img[ 1174] = 238;
assign img[ 1175] = 254;
assign img[ 1176] = 255;
assign img[ 1177] = 255;
assign img[ 1178] = 170;
assign img[ 1179] = 238;
assign img[ 1180] = 238;
assign img[ 1181] = 255;
assign img[ 1182] = 223;
assign img[ 1183] = 157;
assign img[ 1184] = 217;
assign img[ 1185] = 252;
assign img[ 1186] = 238;
assign img[ 1187] = 238;
assign img[ 1188] = 238;
assign img[ 1189] = 239;
assign img[ 1190] = 238;
assign img[ 1191] = 255;
assign img[ 1192] = 255;
assign img[ 1193] = 255;
assign img[ 1194] = 255;
assign img[ 1195] = 255;
assign img[ 1196] = 255;
assign img[ 1197] = 255;
assign img[ 1198] = 255;
assign img[ 1199] = 255;
assign img[ 1200] = 238;
assign img[ 1201] = 238;
assign img[ 1202] = 254;
assign img[ 1203] = 223;
assign img[ 1204] = 204;
assign img[ 1205] = 204;
assign img[ 1206] = 236;
assign img[ 1207] = 255;
assign img[ 1208] = 255;
assign img[ 1209] = 223;
assign img[ 1210] = 239;
assign img[ 1211] = 238;
assign img[ 1212] = 238;
assign img[ 1213] = 207;
assign img[ 1214] = 238;
assign img[ 1215] = 255;
assign img[ 1216] = 255;
assign img[ 1217] = 255;
assign img[ 1218] = 239;
assign img[ 1219] = 238;
assign img[ 1220] = 238;
assign img[ 1221] = 238;
assign img[ 1222] = 238;
assign img[ 1223] = 238;
assign img[ 1224] = 238;
assign img[ 1225] = 238;
assign img[ 1226] = 238;
assign img[ 1227] = 207;
assign img[ 1228] = 204;
assign img[ 1229] = 238;
assign img[ 1230] = 238;
assign img[ 1231] = 238;
assign img[ 1232] = 238;
assign img[ 1233] = 238;
assign img[ 1234] = 206;
assign img[ 1235] = 204;
assign img[ 1236] = 220;
assign img[ 1237] = 205;
assign img[ 1238] = 236;
assign img[ 1239] = 238;
assign img[ 1240] = 238;
assign img[ 1241] = 238;
assign img[ 1242] = 238;
assign img[ 1243] = 254;
assign img[ 1244] = 255;
assign img[ 1245] = 255;
assign img[ 1246] = 238;
assign img[ 1247] = 238;
assign img[ 1248] = 254;
assign img[ 1249] = 255;
assign img[ 1250] = 255;
assign img[ 1251] = 255;
assign img[ 1252] = 255;
assign img[ 1253] = 255;
assign img[ 1254] = 255;
assign img[ 1255] = 255;
assign img[ 1256] = 255;
assign img[ 1257] = 255;
assign img[ 1258] = 255;
assign img[ 1259] = 255;
assign img[ 1260] = 191;
assign img[ 1261] = 255;
assign img[ 1262] = 239;
assign img[ 1263] = 255;
assign img[ 1264] = 239;
assign img[ 1265] = 238;
assign img[ 1266] = 238;
assign img[ 1267] = 255;
assign img[ 1268] = 221;
assign img[ 1269] = 253;
assign img[ 1270] = 255;
assign img[ 1271] = 255;
assign img[ 1272] = 255;
assign img[ 1273] = 191;
assign img[ 1274] = 155;
assign img[ 1275] = 221;
assign img[ 1276] = 205;
assign img[ 1277] = 236;
assign img[ 1278] = 142;
assign img[ 1279] = 236;
assign img[ 1280] = 96;
assign img[ 1281] = 206;
assign img[ 1282] = 236;
assign img[ 1283] = 238;
assign img[ 1284] = 238;
assign img[ 1285] = 254;
assign img[ 1286] = 221;
assign img[ 1287] = 239;
assign img[ 1288] = 238;
assign img[ 1289] = 239;
assign img[ 1290] = 238;
assign img[ 1291] = 238;
assign img[ 1292] = 206;
assign img[ 1293] = 204;
assign img[ 1294] = 220;
assign img[ 1295] = 221;
assign img[ 1296] = 205;
assign img[ 1297] = 220;
assign img[ 1298] = 221;
assign img[ 1299] = 205;
assign img[ 1300] = 236;
assign img[ 1301] = 254;
assign img[ 1302] = 221;
assign img[ 1303] = 253;
assign img[ 1304] = 254;
assign img[ 1305] = 255;
assign img[ 1306] = 255;
assign img[ 1307] = 255;
assign img[ 1308] = 239;
assign img[ 1309] = 255;
assign img[ 1310] = 255;
assign img[ 1311] = 239;
assign img[ 1312] = 153;
assign img[ 1313] = 251;
assign img[ 1314] = 255;
assign img[ 1315] = 255;
assign img[ 1316] = 255;
assign img[ 1317] = 255;
assign img[ 1318] = 255;
assign img[ 1319] = 255;
assign img[ 1320] = 255;
assign img[ 1321] = 255;
assign img[ 1322] = 239;
assign img[ 1323] = 238;
assign img[ 1324] = 254;
assign img[ 1325] = 223;
assign img[ 1326] = 255;
assign img[ 1327] = 207;
assign img[ 1328] = 252;
assign img[ 1329] = 255;
assign img[ 1330] = 239;
assign img[ 1331] = 223;
assign img[ 1332] = 253;
assign img[ 1333] = 255;
assign img[ 1334] = 255;
assign img[ 1335] = 239;
assign img[ 1336] = 238;
assign img[ 1337] = 239;
assign img[ 1338] = 254;
assign img[ 1339] = 255;
assign img[ 1340] = 255;
assign img[ 1341] = 255;
assign img[ 1342] = 255;
assign img[ 1343] = 255;
assign img[ 1344] = 255;
assign img[ 1345] = 255;
assign img[ 1346] = 255;
assign img[ 1347] = 255;
assign img[ 1348] = 255;
assign img[ 1349] = 239;
assign img[ 1350] = 238;
assign img[ 1351] = 238;
assign img[ 1352] = 238;
assign img[ 1353] = 238;
assign img[ 1354] = 254;
assign img[ 1355] = 255;
assign img[ 1356] = 223;
assign img[ 1357] = 221;
assign img[ 1358] = 236;
assign img[ 1359] = 255;
assign img[ 1360] = 255;
assign img[ 1361] = 255;
assign img[ 1362] = 223;
assign img[ 1363] = 255;
assign img[ 1364] = 255;
assign img[ 1365] = 255;
assign img[ 1366] = 238;
assign img[ 1367] = 238;
assign img[ 1368] = 255;
assign img[ 1369] = 255;
assign img[ 1370] = 191;
assign img[ 1371] = 223;
assign img[ 1372] = 253;
assign img[ 1373] = 239;
assign img[ 1374] = 238;
assign img[ 1375] = 174;
assign img[ 1376] = 238;
assign img[ 1377] = 238;
assign img[ 1378] = 254;
assign img[ 1379] = 255;
assign img[ 1380] = 238;
assign img[ 1381] = 255;
assign img[ 1382] = 223;
assign img[ 1383] = 255;
assign img[ 1384] = 255;
assign img[ 1385] = 223;
assign img[ 1386] = 205;
assign img[ 1387] = 204;
assign img[ 1388] = 204;
assign img[ 1389] = 220;
assign img[ 1390] = 221;
assign img[ 1391] = 221;
assign img[ 1392] = 204;
assign img[ 1393] = 206;
assign img[ 1394] = 238;
assign img[ 1395] = 206;
assign img[ 1396] = 204;
assign img[ 1397] = 238;
assign img[ 1398] = 238;
assign img[ 1399] = 254;
assign img[ 1400] = 255;
assign img[ 1401] = 255;
assign img[ 1402] = 223;
assign img[ 1403] = 221;
assign img[ 1404] = 221;
assign img[ 1405] = 253;
assign img[ 1406] = 223;
assign img[ 1407] = 253;
assign img[ 1408] = 96;
assign img[ 1409] = 191;
assign img[ 1410] = 251;
assign img[ 1411] = 255;
assign img[ 1412] = 204;
assign img[ 1413] = 204;
assign img[ 1414] = 204;
assign img[ 1415] = 253;
assign img[ 1416] = 255;
assign img[ 1417] = 255;
assign img[ 1418] = 239;
assign img[ 1419] = 174;
assign img[ 1420] = 170;
assign img[ 1421] = 238;
assign img[ 1422] = 174;
assign img[ 1423] = 206;
assign img[ 1424] = 254;
assign img[ 1425] = 207;
assign img[ 1426] = 220;
assign img[ 1427] = 221;
assign img[ 1428] = 237;
assign img[ 1429] = 238;
assign img[ 1430] = 238;
assign img[ 1431] = 238;
assign img[ 1432] = 254;
assign img[ 1433] = 255;
assign img[ 1434] = 155;
assign img[ 1435] = 255;
assign img[ 1436] = 255;
assign img[ 1437] = 255;
assign img[ 1438] = 223;
assign img[ 1439] = 207;
assign img[ 1440] = 140;
assign img[ 1441] = 238;
assign img[ 1442] = 238;
assign img[ 1443] = 238;
assign img[ 1444] = 254;
assign img[ 1445] = 239;
assign img[ 1446] = 238;
assign img[ 1447] = 255;
assign img[ 1448] = 255;
assign img[ 1449] = 255;
assign img[ 1450] = 255;
assign img[ 1451] = 255;
assign img[ 1452] = 239;
assign img[ 1453] = 238;
assign img[ 1454] = 238;
assign img[ 1455] = 239;
assign img[ 1456] = 255;
assign img[ 1457] = 255;
assign img[ 1458] = 255;
assign img[ 1459] = 255;
assign img[ 1460] = 255;
assign img[ 1461] = 255;
assign img[ 1462] = 238;
assign img[ 1463] = 238;
assign img[ 1464] = 254;
assign img[ 1465] = 255;
assign img[ 1466] = 255;
assign img[ 1467] = 255;
assign img[ 1468] = 255;
assign img[ 1469] = 239;
assign img[ 1470] = 238;
assign img[ 1471] = 255;
assign img[ 1472] = 255;
assign img[ 1473] = 255;
assign img[ 1474] = 239;
assign img[ 1475] = 238;
assign img[ 1476] = 238;
assign img[ 1477] = 206;
assign img[ 1478] = 236;
assign img[ 1479] = 238;
assign img[ 1480] = 238;
assign img[ 1481] = 238;
assign img[ 1482] = 238;
assign img[ 1483] = 238;
assign img[ 1484] = 238;
assign img[ 1485] = 238;
assign img[ 1486] = 238;
assign img[ 1487] = 255;
assign img[ 1488] = 239;
assign img[ 1489] = 238;
assign img[ 1490] = 238;
assign img[ 1491] = 239;
assign img[ 1492] = 223;
assign img[ 1493] = 239;
assign img[ 1494] = 238;
assign img[ 1495] = 238;
assign img[ 1496] = 206;
assign img[ 1497] = 238;
assign img[ 1498] = 238;
assign img[ 1499] = 206;
assign img[ 1500] = 236;
assign img[ 1501] = 238;
assign img[ 1502] = 238;
assign img[ 1503] = 174;
assign img[ 1504] = 136;
assign img[ 1505] = 136;
assign img[ 1506] = 232;
assign img[ 1507] = 255;
assign img[ 1508] = 238;
assign img[ 1509] = 255;
assign img[ 1510] = 204;
assign img[ 1511] = 238;
assign img[ 1512] = 254;
assign img[ 1513] = 255;
assign img[ 1514] = 255;
assign img[ 1515] = 255;
assign img[ 1516] = 206;
assign img[ 1517] = 238;
assign img[ 1518] = 255;
assign img[ 1519] = 207;
assign img[ 1520] = 220;
assign img[ 1521] = 221;
assign img[ 1522] = 221;
assign img[ 1523] = 255;
assign img[ 1524] = 191;
assign img[ 1525] = 187;
assign img[ 1526] = 234;
assign img[ 1527] = 206;
assign img[ 1528] = 220;
assign img[ 1529] = 221;
assign img[ 1530] = 169;
assign img[ 1531] = 238;
assign img[ 1532] = 170;
assign img[ 1533] = 254;
assign img[ 1534] = 191;
assign img[ 1535] = 255;
assign img[ 1536] = 112;
assign img[ 1537] = 239;
assign img[ 1538] = 238;
assign img[ 1539] = 255;
assign img[ 1540] = 255;
assign img[ 1541] = 255;
assign img[ 1542] = 157;
assign img[ 1543] = 255;
assign img[ 1544] = 255;
assign img[ 1545] = 255;
assign img[ 1546] = 255;
assign img[ 1547] = 255;
assign img[ 1548] = 255;
assign img[ 1549] = 255;
assign img[ 1550] = 239;
assign img[ 1551] = 238;
assign img[ 1552] = 238;
assign img[ 1553] = 238;
assign img[ 1554] = 238;
assign img[ 1555] = 255;
assign img[ 1556] = 239;
assign img[ 1557] = 238;
assign img[ 1558] = 238;
assign img[ 1559] = 238;
assign img[ 1560] = 238;
assign img[ 1561] = 238;
assign img[ 1562] = 254;
assign img[ 1563] = 255;
assign img[ 1564] = 255;
assign img[ 1565] = 255;
assign img[ 1566] = 239;
assign img[ 1567] = 255;
assign img[ 1568] = 187;
assign img[ 1569] = 251;
assign img[ 1570] = 207;
assign img[ 1571] = 238;
assign img[ 1572] = 238;
assign img[ 1573] = 206;
assign img[ 1574] = 220;
assign img[ 1575] = 255;
assign img[ 1576] = 255;
assign img[ 1577] = 255;
assign img[ 1578] = 238;
assign img[ 1579] = 238;
assign img[ 1580] = 238;
assign img[ 1581] = 206;
assign img[ 1582] = 236;
assign img[ 1583] = 206;
assign img[ 1584] = 236;
assign img[ 1585] = 255;
assign img[ 1586] = 255;
assign img[ 1587] = 255;
assign img[ 1588] = 255;
assign img[ 1589] = 255;
assign img[ 1590] = 255;
assign img[ 1591] = 255;
assign img[ 1592] = 255;
assign img[ 1593] = 255;
assign img[ 1594] = 255;
assign img[ 1595] = 254;
assign img[ 1596] = 254;
assign img[ 1597] = 255;
assign img[ 1598] = 254;
assign img[ 1599] = 255;
assign img[ 1600] = 255;
assign img[ 1601] = 255;
assign img[ 1602] = 255;
assign img[ 1603] = 255;
assign img[ 1604] = 255;
assign img[ 1605] = 175;
assign img[ 1606] = 186;
assign img[ 1607] = 239;
assign img[ 1608] = 254;
assign img[ 1609] = 255;
assign img[ 1610] = 255;
assign img[ 1611] = 255;
assign img[ 1612] = 255;
assign img[ 1613] = 255;
assign img[ 1614] = 254;
assign img[ 1615] = 254;
assign img[ 1616] = 255;
assign img[ 1617] = 255;
assign img[ 1618] = 255;
assign img[ 1619] = 239;
assign img[ 1620] = 238;
assign img[ 1621] = 238;
assign img[ 1622] = 238;
assign img[ 1623] = 238;
assign img[ 1624] = 254;
assign img[ 1625] = 255;
assign img[ 1626] = 255;
assign img[ 1627] = 255;
assign img[ 1628] = 238;
assign img[ 1629] = 255;
assign img[ 1630] = 255;
assign img[ 1631] = 191;
assign img[ 1632] = 255;
assign img[ 1633] = 255;
assign img[ 1634] = 255;
assign img[ 1635] = 255;
assign img[ 1636] = 255;
assign img[ 1637] = 255;
assign img[ 1638] = 155;
assign img[ 1639] = 255;
assign img[ 1640] = 255;
assign img[ 1641] = 255;
assign img[ 1642] = 238;
assign img[ 1643] = 238;
assign img[ 1644] = 254;
assign img[ 1645] = 255;
assign img[ 1646] = 255;
assign img[ 1647] = 255;
assign img[ 1648] = 255;
assign img[ 1649] = 255;
assign img[ 1650] = 238;
assign img[ 1651] = 238;
assign img[ 1652] = 254;
assign img[ 1653] = 255;
assign img[ 1654] = 255;
assign img[ 1655] = 255;
assign img[ 1656] = 238;
assign img[ 1657] = 255;
assign img[ 1658] = 255;
assign img[ 1659] = 255;
assign img[ 1660] = 255;
assign img[ 1661] = 255;
assign img[ 1662] = 255;
assign img[ 1663] = 255;
assign img[ 1664] = 96;
assign img[ 1665] = 206;
assign img[ 1666] = 236;
assign img[ 1667] = 206;
assign img[ 1668] = 204;
assign img[ 1669] = 221;
assign img[ 1670] = 189;
assign img[ 1671] = 238;
assign img[ 1672] = 238;
assign img[ 1673] = 238;
assign img[ 1674] = 238;
assign img[ 1675] = 255;
assign img[ 1676] = 205;
assign img[ 1677] = 204;
assign img[ 1678] = 236;
assign img[ 1679] = 238;
assign img[ 1680] = 220;
assign img[ 1681] = 239;
assign img[ 1682] = 238;
assign img[ 1683] = 255;
assign img[ 1684] = 255;
assign img[ 1685] = 255;
assign img[ 1686] = 223;
assign img[ 1687] = 255;
assign img[ 1688] = 255;
assign img[ 1689] = 239;
assign img[ 1690] = 238;
assign img[ 1691] = 238;
assign img[ 1692] = 238;
assign img[ 1693] = 238;
assign img[ 1694] = 238;
assign img[ 1695] = 254;
assign img[ 1696] = 187;
assign img[ 1697] = 171;
assign img[ 1698] = 234;
assign img[ 1699] = 255;
assign img[ 1700] = 239;
assign img[ 1701] = 142;
assign img[ 1702] = 232;
assign img[ 1703] = 239;
assign img[ 1704] = 238;
assign img[ 1705] = 238;
assign img[ 1706] = 238;
assign img[ 1707] = 238;
assign img[ 1708] = 238;
assign img[ 1709] = 254;
assign img[ 1710] = 238;
assign img[ 1711] = 255;
assign img[ 1712] = 255;
assign img[ 1713] = 255;
assign img[ 1714] = 255;
assign img[ 1715] = 255;
assign img[ 1716] = 239;
assign img[ 1717] = 238;
assign img[ 1718] = 238;
assign img[ 1719] = 238;
assign img[ 1720] = 254;
assign img[ 1721] = 255;
assign img[ 1722] = 239;
assign img[ 1723] = 238;
assign img[ 1724] = 238;
assign img[ 1725] = 239;
assign img[ 1726] = 238;
assign img[ 1727] = 255;
assign img[ 1728] = 255;
assign img[ 1729] = 255;
assign img[ 1730] = 239;
assign img[ 1731] = 238;
assign img[ 1732] = 238;
assign img[ 1733] = 238;
assign img[ 1734] = 220;
assign img[ 1735] = 221;
assign img[ 1736] = 221;
assign img[ 1737] = 255;
assign img[ 1738] = 255;
assign img[ 1739] = 255;
assign img[ 1740] = 238;
assign img[ 1741] = 255;
assign img[ 1742] = 255;
assign img[ 1743] = 255;
assign img[ 1744] = 255;
assign img[ 1745] = 255;
assign img[ 1746] = 223;
assign img[ 1747] = 255;
assign img[ 1748] = 255;
assign img[ 1749] = 255;
assign img[ 1750] = 255;
assign img[ 1751] = 255;
assign img[ 1752] = 239;
assign img[ 1753] = 255;
assign img[ 1754] = 175;
assign img[ 1755] = 238;
assign img[ 1756] = 238;
assign img[ 1757] = 238;
assign img[ 1758] = 238;
assign img[ 1759] = 191;
assign img[ 1760] = 187;
assign img[ 1761] = 255;
assign img[ 1762] = 255;
assign img[ 1763] = 255;
assign img[ 1764] = 255;
assign img[ 1765] = 255;
assign img[ 1766] = 223;
assign img[ 1767] = 255;
assign img[ 1768] = 255;
assign img[ 1769] = 255;
assign img[ 1770] = 255;
assign img[ 1771] = 255;
assign img[ 1772] = 255;
assign img[ 1773] = 255;
assign img[ 1774] = 255;
assign img[ 1775] = 255;
assign img[ 1776] = 239;
assign img[ 1777] = 255;
assign img[ 1778] = 239;
assign img[ 1779] = 238;
assign img[ 1780] = 238;
assign img[ 1781] = 238;
assign img[ 1782] = 238;
assign img[ 1783] = 238;
assign img[ 1784] = 238;
assign img[ 1785] = 174;
assign img[ 1786] = 170;
assign img[ 1787] = 138;
assign img[ 1788] = 200;
assign img[ 1789] = 236;
assign img[ 1790] = 222;
assign img[ 1791] = 253;
assign img[ 1792] = 96;
assign img[ 1793] = 206;
assign img[ 1794] = 236;
assign img[ 1795] = 238;
assign img[ 1796] = 254;
assign img[ 1797] = 223;
assign img[ 1798] = 221;
assign img[ 1799] = 255;
assign img[ 1800] = 255;
assign img[ 1801] = 255;
assign img[ 1802] = 239;
assign img[ 1803] = 254;
assign img[ 1804] = 239;
assign img[ 1805] = 238;
assign img[ 1806] = 238;
assign img[ 1807] = 206;
assign img[ 1808] = 204;
assign img[ 1809] = 204;
assign img[ 1810] = 236;
assign img[ 1811] = 238;
assign img[ 1812] = 238;
assign img[ 1813] = 254;
assign img[ 1814] = 221;
assign img[ 1815] = 253;
assign img[ 1816] = 255;
assign img[ 1817] = 255;
assign img[ 1818] = 239;
assign img[ 1819] = 238;
assign img[ 1820] = 238;
assign img[ 1821] = 238;
assign img[ 1822] = 238;
assign img[ 1823] = 238;
assign img[ 1824] = 220;
assign img[ 1825] = 253;
assign img[ 1826] = 255;
assign img[ 1827] = 255;
assign img[ 1828] = 239;
assign img[ 1829] = 255;
assign img[ 1830] = 255;
assign img[ 1831] = 206;
assign img[ 1832] = 236;
assign img[ 1833] = 255;
assign img[ 1834] = 255;
assign img[ 1835] = 255;
assign img[ 1836] = 255;
assign img[ 1837] = 255;
assign img[ 1838] = 238;
assign img[ 1839] = 255;
assign img[ 1840] = 255;
assign img[ 1841] = 255;
assign img[ 1842] = 255;
assign img[ 1843] = 255;
assign img[ 1844] = 255;
assign img[ 1845] = 255;
assign img[ 1846] = 255;
assign img[ 1847] = 255;
assign img[ 1848] = 255;
assign img[ 1849] = 255;
assign img[ 1850] = 255;
assign img[ 1851] = 255;
assign img[ 1852] = 255;
assign img[ 1853] = 223;
assign img[ 1854] = 255;
assign img[ 1855] = 255;
assign img[ 1856] = 255;
assign img[ 1857] = 255;
assign img[ 1858] = 255;
assign img[ 1859] = 255;
assign img[ 1860] = 255;
assign img[ 1861] = 239;
assign img[ 1862] = 238;
assign img[ 1863] = 255;
assign img[ 1864] = 255;
assign img[ 1865] = 255;
assign img[ 1866] = 255;
assign img[ 1867] = 255;
assign img[ 1868] = 255;
assign img[ 1869] = 255;
assign img[ 1870] = 255;
assign img[ 1871] = 255;
assign img[ 1872] = 255;
assign img[ 1873] = 255;
assign img[ 1874] = 255;
assign img[ 1875] = 255;
assign img[ 1876] = 255;
assign img[ 1877] = 255;
assign img[ 1878] = 255;
assign img[ 1879] = 255;
assign img[ 1880] = 255;
assign img[ 1881] = 239;
assign img[ 1882] = 238;
assign img[ 1883] = 238;
assign img[ 1884] = 238;
assign img[ 1885] = 238;
assign img[ 1886] = 238;
assign img[ 1887] = 238;
assign img[ 1888] = 255;
assign img[ 1889] = 238;
assign img[ 1890] = 238;
assign img[ 1891] = 238;
assign img[ 1892] = 238;
assign img[ 1893] = 255;
assign img[ 1894] = 255;
assign img[ 1895] = 255;
assign img[ 1896] = 255;
assign img[ 1897] = 255;
assign img[ 1898] = 255;
assign img[ 1899] = 255;
assign img[ 1900] = 191;
assign img[ 1901] = 255;
assign img[ 1902] = 255;
assign img[ 1903] = 255;
assign img[ 1904] = 239;
assign img[ 1905] = 239;
assign img[ 1906] = 238;
assign img[ 1907] = 239;
assign img[ 1908] = 255;
assign img[ 1909] = 255;
assign img[ 1910] = 238;
assign img[ 1911] = 238;
assign img[ 1912] = 254;
assign img[ 1913] = 255;
assign img[ 1914] = 255;
assign img[ 1915] = 255;
assign img[ 1916] = 221;
assign img[ 1917] = 255;
assign img[ 1918] = 223;
assign img[ 1919] = 255;
assign img[ 1920] = 96;
assign img[ 1921] = 239;
assign img[ 1922] = 238;
assign img[ 1923] = 238;
assign img[ 1924] = 222;
assign img[ 1925] = 223;
assign img[ 1926] = 221;
assign img[ 1927] = 255;
assign img[ 1928] = 255;
assign img[ 1929] = 255;
assign img[ 1930] = 255;
assign img[ 1931] = 191;
assign img[ 1932] = 155;
assign img[ 1933] = 187;
assign img[ 1934] = 187;
assign img[ 1935] = 223;
assign img[ 1936] = 221;
assign img[ 1937] = 221;
assign img[ 1938] = 236;
assign img[ 1939] = 255;
assign img[ 1940] = 187;
assign img[ 1941] = 255;
assign img[ 1942] = 255;
assign img[ 1943] = 255;
assign img[ 1944] = 255;
assign img[ 1945] = 239;
assign img[ 1946] = 238;
assign img[ 1947] = 238;
assign img[ 1948] = 204;
assign img[ 1949] = 254;
assign img[ 1950] = 223;
assign img[ 1951] = 205;
assign img[ 1952] = 204;
assign img[ 1953] = 253;
assign img[ 1954] = 255;
assign img[ 1955] = 255;
assign img[ 1956] = 239;
assign img[ 1957] = 238;
assign img[ 1958] = 254;
assign img[ 1959] = 255;
assign img[ 1960] = 238;
assign img[ 1961] = 255;
assign img[ 1962] = 255;
assign img[ 1963] = 255;
assign img[ 1964] = 255;
assign img[ 1965] = 223;
assign img[ 1966] = 253;
assign img[ 1967] = 223;
assign img[ 1968] = 253;
assign img[ 1969] = 255;
assign img[ 1970] = 255;
assign img[ 1971] = 255;
assign img[ 1972] = 255;
assign img[ 1973] = 255;
assign img[ 1974] = 255;
assign img[ 1975] = 255;
assign img[ 1976] = 255;
assign img[ 1977] = 255;
assign img[ 1978] = 239;
assign img[ 1979] = 238;
assign img[ 1980] = 238;
assign img[ 1981] = 238;
assign img[ 1982] = 238;
assign img[ 1983] = 255;
assign img[ 1984] = 255;
assign img[ 1985] = 255;
assign img[ 1986] = 255;
assign img[ 1987] = 255;
assign img[ 1988] = 255;
assign img[ 1989] = 255;
assign img[ 1990] = 255;
assign img[ 1991] = 255;
assign img[ 1992] = 255;
assign img[ 1993] = 255;
assign img[ 1994] = 255;
assign img[ 1995] = 255;
assign img[ 1996] = 221;
assign img[ 1997] = 239;
assign img[ 1998] = 238;
assign img[ 1999] = 255;
assign img[ 2000] = 223;
assign img[ 2001] = 255;
assign img[ 2002] = 255;
assign img[ 2003] = 255;
assign img[ 2004] = 205;
assign img[ 2005] = 204;
assign img[ 2006] = 204;
assign img[ 2007] = 236;
assign img[ 2008] = 206;
assign img[ 2009] = 236;
assign img[ 2010] = 254;
assign img[ 2011] = 255;
assign img[ 2012] = 255;
assign img[ 2013] = 255;
assign img[ 2014] = 255;
assign img[ 2015] = 255;
assign img[ 2016] = 153;
assign img[ 2017] = 137;
assign img[ 2018] = 253;
assign img[ 2019] = 255;
assign img[ 2020] = 239;
assign img[ 2021] = 239;
assign img[ 2022] = 255;
assign img[ 2023] = 255;
assign img[ 2024] = 255;
assign img[ 2025] = 255;
assign img[ 2026] = 255;
assign img[ 2027] = 255;
assign img[ 2028] = 255;
assign img[ 2029] = 255;
assign img[ 2030] = 239;
assign img[ 2031] = 238;
assign img[ 2032] = 204;
assign img[ 2033] = 236;
assign img[ 2034] = 170;
assign img[ 2035] = 187;
assign img[ 2036] = 187;
assign img[ 2037] = 187;
assign img[ 2038] = 251;
assign img[ 2039] = 255;
assign img[ 2040] = 255;
assign img[ 2041] = 255;
assign img[ 2042] = 155;
assign img[ 2043] = 153;
assign img[ 2044] = 221;
assign img[ 2045] = 255;
assign img[ 2046] = 239;
assign img[ 2047] = 238;
assign img[ 2048] = 96;
assign img[ 2049] = 238;
assign img[ 2050] = 254;
assign img[ 2051] = 239;
assign img[ 2052] = 174;
assign img[ 2053] = 254;
assign img[ 2054] = 159;
assign img[ 2055] = 255;
assign img[ 2056] = 255;
assign img[ 2057] = 255;
assign img[ 2058] = 255;
assign img[ 2059] = 223;
assign img[ 2060] = 205;
assign img[ 2061] = 204;
assign img[ 2062] = 236;
assign img[ 2063] = 206;
assign img[ 2064] = 236;
assign img[ 2065] = 206;
assign img[ 2066] = 236;
assign img[ 2067] = 255;
assign img[ 2068] = 139;
assign img[ 2069] = 238;
assign img[ 2070] = 238;
assign img[ 2071] = 254;
assign img[ 2072] = 255;
assign img[ 2073] = 255;
assign img[ 2074] = 187;
assign img[ 2075] = 255;
assign img[ 2076] = 255;
assign img[ 2077] = 255;
assign img[ 2078] = 255;
assign img[ 2079] = 255;
assign img[ 2080] = 103;
assign img[ 2081] = 230;
assign img[ 2082] = 238;
assign img[ 2083] = 238;
assign img[ 2084] = 206;
assign img[ 2085] = 238;
assign img[ 2086] = 238;
assign img[ 2087] = 238;
assign img[ 2088] = 238;
assign img[ 2089] = 238;
assign img[ 2090] = 190;
assign img[ 2091] = 171;
assign img[ 2092] = 234;
assign img[ 2093] = 238;
assign img[ 2094] = 238;
assign img[ 2095] = 238;
assign img[ 2096] = 238;
assign img[ 2097] = 238;
assign img[ 2098] = 238;
assign img[ 2099] = 238;
assign img[ 2100] = 206;
assign img[ 2101] = 238;
assign img[ 2102] = 238;
assign img[ 2103] = 207;
assign img[ 2104] = 252;
assign img[ 2105] = 255;
assign img[ 2106] = 238;
assign img[ 2107] = 238;
assign img[ 2108] = 238;
assign img[ 2109] = 255;
assign img[ 2110] = 255;
assign img[ 2111] = 255;
assign img[ 2112] = 255;
assign img[ 2113] = 255;
assign img[ 2114] = 191;
assign img[ 2115] = 255;
assign img[ 2116] = 255;
assign img[ 2117] = 255;
assign img[ 2118] = 238;
assign img[ 2119] = 238;
assign img[ 2120] = 255;
assign img[ 2121] = 255;
assign img[ 2122] = 255;
assign img[ 2123] = 255;
assign img[ 2124] = 255;
assign img[ 2125] = 255;
assign img[ 2126] = 255;
assign img[ 2127] = 255;
assign img[ 2128] = 255;
assign img[ 2129] = 255;
assign img[ 2130] = 255;
assign img[ 2131] = 255;
assign img[ 2132] = 255;
assign img[ 2133] = 191;
assign img[ 2134] = 251;
assign img[ 2135] = 255;
assign img[ 2136] = 255;
assign img[ 2137] = 255;
assign img[ 2138] = 255;
assign img[ 2139] = 255;
assign img[ 2140] = 255;
assign img[ 2141] = 255;
assign img[ 2142] = 255;
assign img[ 2143] = 255;
assign img[ 2144] = 187;
assign img[ 2145] = 119;
assign img[ 2146] = 247;
assign img[ 2147] = 255;
assign img[ 2148] = 255;
assign img[ 2149] = 239;
assign img[ 2150] = 238;
assign img[ 2151] = 238;
assign img[ 2152] = 254;
assign img[ 2153] = 239;
assign img[ 2154] = 238;
assign img[ 2155] = 238;
assign img[ 2156] = 238;
assign img[ 2157] = 238;
assign img[ 2158] = 238;
assign img[ 2159] = 238;
assign img[ 2160] = 223;
assign img[ 2161] = 205;
assign img[ 2162] = 236;
assign img[ 2163] = 206;
assign img[ 2164] = 204;
assign img[ 2165] = 204;
assign img[ 2166] = 236;
assign img[ 2167] = 238;
assign img[ 2168] = 238;
assign img[ 2169] = 239;
assign img[ 2170] = 238;
assign img[ 2171] = 191;
assign img[ 2172] = 255;
assign img[ 2173] = 255;
assign img[ 2174] = 255;
assign img[ 2175] = 255;
assign img[ 2176] = 96;
assign img[ 2177] = 239;
assign img[ 2178] = 238;
assign img[ 2179] = 238;
assign img[ 2180] = 254;
assign img[ 2181] = 255;
assign img[ 2182] = 207;
assign img[ 2183] = 238;
assign img[ 2184] = 238;
assign img[ 2185] = 238;
assign img[ 2186] = 238;
assign img[ 2187] = 238;
assign img[ 2188] = 206;
assign img[ 2189] = 238;
assign img[ 2190] = 158;
assign img[ 2191] = 221;
assign img[ 2192] = 236;
assign img[ 2193] = 255;
assign img[ 2194] = 255;
assign img[ 2195] = 239;
assign img[ 2196] = 254;
assign img[ 2197] = 255;
assign img[ 2198] = 255;
assign img[ 2199] = 255;
assign img[ 2200] = 255;
assign img[ 2201] = 255;
assign img[ 2202] = 238;
assign img[ 2203] = 238;
assign img[ 2204] = 238;
assign img[ 2205] = 254;
assign img[ 2206] = 239;
assign img[ 2207] = 191;
assign img[ 2208] = 187;
assign img[ 2209] = 234;
assign img[ 2210] = 238;
assign img[ 2211] = 238;
assign img[ 2212] = 238;
assign img[ 2213] = 238;
assign img[ 2214] = 238;
assign img[ 2215] = 254;
assign img[ 2216] = 255;
assign img[ 2217] = 255;
assign img[ 2218] = 142;
assign img[ 2219] = 238;
assign img[ 2220] = 238;
assign img[ 2221] = 238;
assign img[ 2222] = 238;
assign img[ 2223] = 238;
assign img[ 2224] = 254;
assign img[ 2225] = 255;
assign img[ 2226] = 255;
assign img[ 2227] = 255;
assign img[ 2228] = 255;
assign img[ 2229] = 255;
assign img[ 2230] = 255;
assign img[ 2231] = 255;
assign img[ 2232] = 239;
assign img[ 2233] = 238;
assign img[ 2234] = 238;
assign img[ 2235] = 238;
assign img[ 2236] = 238;
assign img[ 2237] = 255;
assign img[ 2238] = 255;
assign img[ 2239] = 255;
assign img[ 2240] = 255;
assign img[ 2241] = 239;
assign img[ 2242] = 238;
assign img[ 2243] = 238;
assign img[ 2244] = 238;
assign img[ 2245] = 238;
assign img[ 2246] = 238;
assign img[ 2247] = 238;
assign img[ 2248] = 238;
assign img[ 2249] = 238;
assign img[ 2250] = 238;
assign img[ 2251] = 255;
assign img[ 2252] = 255;
assign img[ 2253] = 255;
assign img[ 2254] = 255;
assign img[ 2255] = 255;
assign img[ 2256] = 255;
assign img[ 2257] = 255;
assign img[ 2258] = 255;
assign img[ 2259] = 239;
assign img[ 2260] = 238;
assign img[ 2261] = 143;
assign img[ 2262] = 236;
assign img[ 2263] = 238;
assign img[ 2264] = 238;
assign img[ 2265] = 255;
assign img[ 2266] = 238;
assign img[ 2267] = 239;
assign img[ 2268] = 222;
assign img[ 2269] = 254;
assign img[ 2270] = 238;
assign img[ 2271] = 174;
assign img[ 2272] = 186;
assign img[ 2273] = 251;
assign img[ 2274] = 255;
assign img[ 2275] = 255;
assign img[ 2276] = 238;
assign img[ 2277] = 255;
assign img[ 2278] = 255;
assign img[ 2279] = 255;
assign img[ 2280] = 255;
assign img[ 2281] = 255;
assign img[ 2282] = 255;
assign img[ 2283] = 255;
assign img[ 2284] = 255;
assign img[ 2285] = 255;
assign img[ 2286] = 255;
assign img[ 2287] = 255;
assign img[ 2288] = 207;
assign img[ 2289] = 206;
assign img[ 2290] = 238;
assign img[ 2291] = 254;
assign img[ 2292] = 255;
assign img[ 2293] = 255;
assign img[ 2294] = 221;
assign img[ 2295] = 255;
assign img[ 2296] = 255;
assign img[ 2297] = 255;
assign img[ 2298] = 238;
assign img[ 2299] = 238;
assign img[ 2300] = 238;
assign img[ 2301] = 255;
assign img[ 2302] = 238;
assign img[ 2303] = 255;
assign img[ 2304] = 96;
assign img[ 2305] = 238;
assign img[ 2306] = 238;
assign img[ 2307] = 238;
assign img[ 2308] = 252;
assign img[ 2309] = 255;
assign img[ 2310] = 239;
assign img[ 2311] = 254;
assign img[ 2312] = 255;
assign img[ 2313] = 255;
assign img[ 2314] = 255;
assign img[ 2315] = 255;
assign img[ 2316] = 255;
assign img[ 2317] = 255;
assign img[ 2318] = 255;
assign img[ 2319] = 255;
assign img[ 2320] = 187;
assign img[ 2321] = 255;
assign img[ 2322] = 255;
assign img[ 2323] = 255;
assign img[ 2324] = 255;
assign img[ 2325] = 255;
assign img[ 2326] = 255;
assign img[ 2327] = 255;
assign img[ 2328] = 255;
assign img[ 2329] = 239;
assign img[ 2330] = 238;
assign img[ 2331] = 238;
assign img[ 2332] = 238;
assign img[ 2333] = 255;
assign img[ 2334] = 239;
assign img[ 2335] = 206;
assign img[ 2336] = 254;
assign img[ 2337] = 255;
assign img[ 2338] = 254;
assign img[ 2339] = 255;
assign img[ 2340] = 255;
assign img[ 2341] = 255;
assign img[ 2342] = 206;
assign img[ 2343] = 223;
assign img[ 2344] = 255;
assign img[ 2345] = 255;
assign img[ 2346] = 255;
assign img[ 2347] = 255;
assign img[ 2348] = 223;
assign img[ 2349] = 221;
assign img[ 2350] = 236;
assign img[ 2351] = 238;
assign img[ 2352] = 238;
assign img[ 2353] = 255;
assign img[ 2354] = 239;
assign img[ 2355] = 254;
assign img[ 2356] = 255;
assign img[ 2357] = 255;
assign img[ 2358] = 255;
assign img[ 2359] = 255;
assign img[ 2360] = 255;
assign img[ 2361] = 255;
assign img[ 2362] = 255;
assign img[ 2363] = 255;
assign img[ 2364] = 255;
assign img[ 2365] = 255;
assign img[ 2366] = 255;
assign img[ 2367] = 255;
assign img[ 2368] = 255;
assign img[ 2369] = 255;
assign img[ 2370] = 255;
assign img[ 2371] = 255;
assign img[ 2372] = 255;
assign img[ 2373] = 255;
assign img[ 2374] = 221;
assign img[ 2375] = 255;
assign img[ 2376] = 255;
assign img[ 2377] = 255;
assign img[ 2378] = 255;
assign img[ 2379] = 255;
assign img[ 2380] = 255;
assign img[ 2381] = 255;
assign img[ 2382] = 238;
assign img[ 2383] = 238;
assign img[ 2384] = 255;
assign img[ 2385] = 255;
assign img[ 2386] = 238;
assign img[ 2387] = 206;
assign img[ 2388] = 204;
assign img[ 2389] = 206;
assign img[ 2390] = 238;
assign img[ 2391] = 238;
assign img[ 2392] = 238;
assign img[ 2393] = 223;
assign img[ 2394] = 205;
assign img[ 2395] = 204;
assign img[ 2396] = 254;
assign img[ 2397] = 255;
assign img[ 2398] = 255;
assign img[ 2399] = 191;
assign img[ 2400] = 255;
assign img[ 2401] = 255;
assign img[ 2402] = 255;
assign img[ 2403] = 255;
assign img[ 2404] = 255;
assign img[ 2405] = 239;
assign img[ 2406] = 254;
assign img[ 2407] = 238;
assign img[ 2408] = 238;
assign img[ 2409] = 238;
assign img[ 2410] = 238;
assign img[ 2411] = 255;
assign img[ 2412] = 191;
assign img[ 2413] = 255;
assign img[ 2414] = 223;
assign img[ 2415] = 221;
assign img[ 2416] = 255;
assign img[ 2417] = 239;
assign img[ 2418] = 254;
assign img[ 2419] = 255;
assign img[ 2420] = 238;
assign img[ 2421] = 238;
assign img[ 2422] = 238;
assign img[ 2423] = 238;
assign img[ 2424] = 238;
assign img[ 2425] = 255;
assign img[ 2426] = 238;
assign img[ 2427] = 238;
assign img[ 2428] = 254;
assign img[ 2429] = 255;
assign img[ 2430] = 255;
assign img[ 2431] = 255;
assign img[ 2432] = 96;
assign img[ 2433] = 102;
assign img[ 2434] = 118;
assign img[ 2435] = 255;
assign img[ 2436] = 255;
assign img[ 2437] = 255;
assign img[ 2438] = 191;
assign img[ 2439] = 187;
assign img[ 2440] = 234;
assign img[ 2441] = 254;
assign img[ 2442] = 255;
assign img[ 2443] = 255;
assign img[ 2444] = 221;
assign img[ 2445] = 255;
assign img[ 2446] = 255;
assign img[ 2447] = 255;
assign img[ 2448] = 204;
assign img[ 2449] = 238;
assign img[ 2450] = 238;
assign img[ 2451] = 239;
assign img[ 2452] = 204;
assign img[ 2453] = 238;
assign img[ 2454] = 254;
assign img[ 2455] = 255;
assign img[ 2456] = 255;
assign img[ 2457] = 255;
assign img[ 2458] = 238;
assign img[ 2459] = 238;
assign img[ 2460] = 238;
assign img[ 2461] = 255;
assign img[ 2462] = 239;
assign img[ 2463] = 255;
assign img[ 2464] = 187;
assign img[ 2465] = 251;
assign img[ 2466] = 255;
assign img[ 2467] = 255;
assign img[ 2468] = 255;
assign img[ 2469] = 255;
assign img[ 2470] = 255;
assign img[ 2471] = 255;
assign img[ 2472] = 238;
assign img[ 2473] = 238;
assign img[ 2474] = 238;
assign img[ 2475] = 255;
assign img[ 2476] = 255;
assign img[ 2477] = 255;
assign img[ 2478] = 255;
assign img[ 2479] = 223;
assign img[ 2480] = 253;
assign img[ 2481] = 255;
assign img[ 2482] = 255;
assign img[ 2483] = 255;
assign img[ 2484] = 238;
assign img[ 2485] = 238;
assign img[ 2486] = 238;
assign img[ 2487] = 238;
assign img[ 2488] = 238;
assign img[ 2489] = 174;
assign img[ 2490] = 170;
assign img[ 2491] = 255;
assign img[ 2492] = 255;
assign img[ 2493] = 255;
assign img[ 2494] = 221;
assign img[ 2495] = 255;
assign img[ 2496] = 255;
assign img[ 2497] = 255;
assign img[ 2498] = 206;
assign img[ 2499] = 238;
assign img[ 2500] = 254;
assign img[ 2501] = 255;
assign img[ 2502] = 191;
assign img[ 2503] = 187;
assign img[ 2504] = 251;
assign img[ 2505] = 255;
assign img[ 2506] = 255;
assign img[ 2507] = 255;
assign img[ 2508] = 255;
assign img[ 2509] = 255;
assign img[ 2510] = 255;
assign img[ 2511] = 255;
assign img[ 2512] = 223;
assign img[ 2513] = 255;
assign img[ 2514] = 223;
assign img[ 2515] = 205;
assign img[ 2516] = 156;
assign img[ 2517] = 221;
assign img[ 2518] = 253;
assign img[ 2519] = 255;
assign img[ 2520] = 207;
assign img[ 2521] = 238;
assign img[ 2522] = 238;
assign img[ 2523] = 238;
assign img[ 2524] = 238;
assign img[ 2525] = 239;
assign img[ 2526] = 255;
assign img[ 2527] = 255;
assign img[ 2528] = 223;
assign img[ 2529] = 221;
assign img[ 2530] = 253;
assign img[ 2531] = 255;
assign img[ 2532] = 255;
assign img[ 2533] = 255;
assign img[ 2534] = 207;
assign img[ 2535] = 238;
assign img[ 2536] = 254;
assign img[ 2537] = 255;
assign img[ 2538] = 255;
assign img[ 2539] = 255;
assign img[ 2540] = 238;
assign img[ 2541] = 238;
assign img[ 2542] = 238;
assign img[ 2543] = 238;
assign img[ 2544] = 238;
assign img[ 2545] = 238;
assign img[ 2546] = 238;
assign img[ 2547] = 255;
assign img[ 2548] = 255;
assign img[ 2549] = 255;
assign img[ 2550] = 255;
assign img[ 2551] = 255;
assign img[ 2552] = 238;
assign img[ 2553] = 238;
assign img[ 2554] = 238;
assign img[ 2555] = 238;
assign img[ 2556] = 254;
assign img[ 2557] = 255;
assign img[ 2558] = 255;
assign img[ 2559] = 255;
assign img[ 2560] = 96;
assign img[ 2561] = 238;
assign img[ 2562] = 238;
assign img[ 2563] = 223;
assign img[ 2564] = 205;
assign img[ 2565] = 204;
assign img[ 2566] = 204;
assign img[ 2567] = 236;
assign img[ 2568] = 238;
assign img[ 2569] = 255;
assign img[ 2570] = 255;
assign img[ 2571] = 255;
assign img[ 2572] = 255;
assign img[ 2573] = 238;
assign img[ 2574] = 206;
assign img[ 2575] = 204;
assign img[ 2576] = 236;
assign img[ 2577] = 254;
assign img[ 2578] = 255;
assign img[ 2579] = 255;
assign img[ 2580] = 238;
assign img[ 2581] = 238;
assign img[ 2582] = 238;
assign img[ 2583] = 238;
assign img[ 2584] = 238;
assign img[ 2585] = 255;
assign img[ 2586] = 255;
assign img[ 2587] = 255;
assign img[ 2588] = 255;
assign img[ 2589] = 255;
assign img[ 2590] = 255;
assign img[ 2591] = 239;
assign img[ 2592] = 204;
assign img[ 2593] = 254;
assign img[ 2594] = 255;
assign img[ 2595] = 255;
assign img[ 2596] = 238;
assign img[ 2597] = 238;
assign img[ 2598] = 238;
assign img[ 2599] = 238;
assign img[ 2600] = 238;
assign img[ 2601] = 238;
assign img[ 2602] = 238;
assign img[ 2603] = 238;
assign img[ 2604] = 238;
assign img[ 2605] = 239;
assign img[ 2606] = 238;
assign img[ 2607] = 255;
assign img[ 2608] = 255;
assign img[ 2609] = 255;
assign img[ 2610] = 255;
assign img[ 2611] = 255;
assign img[ 2612] = 239;
assign img[ 2613] = 238;
assign img[ 2614] = 238;
assign img[ 2615] = 238;
assign img[ 2616] = 238;
assign img[ 2617] = 254;
assign img[ 2618] = 255;
assign img[ 2619] = 255;
assign img[ 2620] = 255;
assign img[ 2621] = 255;
assign img[ 2622] = 255;
assign img[ 2623] = 255;
assign img[ 2624] = 255;
assign img[ 2625] = 255;
assign img[ 2626] = 223;
assign img[ 2627] = 205;
assign img[ 2628] = 236;
assign img[ 2629] = 238;
assign img[ 2630] = 254;
assign img[ 2631] = 255;
assign img[ 2632] = 255;
assign img[ 2633] = 255;
assign img[ 2634] = 255;
assign img[ 2635] = 239;
assign img[ 2636] = 238;
assign img[ 2637] = 238;
assign img[ 2638] = 238;
assign img[ 2639] = 255;
assign img[ 2640] = 255;
assign img[ 2641] = 255;
assign img[ 2642] = 239;
assign img[ 2643] = 238;
assign img[ 2644] = 238;
assign img[ 2645] = 254;
assign img[ 2646] = 255;
assign img[ 2647] = 255;
assign img[ 2648] = 238;
assign img[ 2649] = 238;
assign img[ 2650] = 238;
assign img[ 2651] = 255;
assign img[ 2652] = 239;
assign img[ 2653] = 238;
assign img[ 2654] = 254;
assign img[ 2655] = 191;
assign img[ 2656] = 255;
assign img[ 2657] = 255;
assign img[ 2658] = 255;
assign img[ 2659] = 255;
assign img[ 2660] = 254;
assign img[ 2661] = 255;
assign img[ 2662] = 254;
assign img[ 2663] = 255;
assign img[ 2664] = 254;
assign img[ 2665] = 255;
assign img[ 2666] = 255;
assign img[ 2667] = 255;
assign img[ 2668] = 255;
assign img[ 2669] = 255;
assign img[ 2670] = 255;
assign img[ 2671] = 255;
assign img[ 2672] = 255;
assign img[ 2673] = 255;
assign img[ 2674] = 221;
assign img[ 2675] = 221;
assign img[ 2676] = 221;
assign img[ 2677] = 221;
assign img[ 2678] = 221;
assign img[ 2679] = 253;
assign img[ 2680] = 239;
assign img[ 2681] = 238;
assign img[ 2682] = 238;
assign img[ 2683] = 254;
assign img[ 2684] = 239;
assign img[ 2685] = 239;
assign img[ 2686] = 255;
assign img[ 2687] = 255;
assign img[ 2688] = 96;
assign img[ 2689] = 239;
assign img[ 2690] = 238;
assign img[ 2691] = 239;
assign img[ 2692] = 221;
assign img[ 2693] = 255;
assign img[ 2694] = 191;
assign img[ 2695] = 255;
assign img[ 2696] = 255;
assign img[ 2697] = 255;
assign img[ 2698] = 255;
assign img[ 2699] = 207;
assign img[ 2700] = 204;
assign img[ 2701] = 204;
assign img[ 2702] = 204;
assign img[ 2703] = 204;
assign img[ 2704] = 156;
assign img[ 2705] = 221;
assign img[ 2706] = 253;
assign img[ 2707] = 255;
assign img[ 2708] = 255;
assign img[ 2709] = 255;
assign img[ 2710] = 255;
assign img[ 2711] = 255;
assign img[ 2712] = 255;
assign img[ 2713] = 191;
assign img[ 2714] = 187;
assign img[ 2715] = 255;
assign img[ 2716] = 255;
assign img[ 2717] = 255;
assign img[ 2718] = 239;
assign img[ 2719] = 174;
assign img[ 2720] = 170;
assign img[ 2721] = 234;
assign img[ 2722] = 238;
assign img[ 2723] = 238;
assign img[ 2724] = 238;
assign img[ 2725] = 238;
assign img[ 2726] = 254;
assign img[ 2727] = 255;
assign img[ 2728] = 255;
assign img[ 2729] = 255;
assign img[ 2730] = 239;
assign img[ 2731] = 238;
assign img[ 2732] = 238;
assign img[ 2733] = 207;
assign img[ 2734] = 238;
assign img[ 2735] = 239;
assign img[ 2736] = 255;
assign img[ 2737] = 255;
assign img[ 2738] = 255;
assign img[ 2739] = 255;
assign img[ 2740] = 239;
assign img[ 2741] = 238;
assign img[ 2742] = 238;
assign img[ 2743] = 238;
assign img[ 2744] = 238;
assign img[ 2745] = 238;
assign img[ 2746] = 254;
assign img[ 2747] = 255;
assign img[ 2748] = 255;
assign img[ 2749] = 239;
assign img[ 2750] = 238;
assign img[ 2751] = 255;
assign img[ 2752] = 255;
assign img[ 2753] = 255;
assign img[ 2754] = 255;
assign img[ 2755] = 255;
assign img[ 2756] = 255;
assign img[ 2757] = 255;
assign img[ 2758] = 255;
assign img[ 2759] = 255;
assign img[ 2760] = 255;
assign img[ 2761] = 255;
assign img[ 2762] = 255;
assign img[ 2763] = 239;
assign img[ 2764] = 238;
assign img[ 2765] = 255;
assign img[ 2766] = 255;
assign img[ 2767] = 255;
assign img[ 2768] = 239;
assign img[ 2769] = 238;
assign img[ 2770] = 206;
assign img[ 2771] = 238;
assign img[ 2772] = 254;
assign img[ 2773] = 255;
assign img[ 2774] = 238;
assign img[ 2775] = 238;
assign img[ 2776] = 238;
assign img[ 2777] = 255;
assign img[ 2778] = 255;
assign img[ 2779] = 255;
assign img[ 2780] = 255;
assign img[ 2781] = 255;
assign img[ 2782] = 255;
assign img[ 2783] = 191;
assign img[ 2784] = 255;
assign img[ 2785] = 251;
assign img[ 2786] = 255;
assign img[ 2787] = 255;
assign img[ 2788] = 255;
assign img[ 2789] = 239;
assign img[ 2790] = 174;
assign img[ 2791] = 238;
assign img[ 2792] = 238;
assign img[ 2793] = 238;
assign img[ 2794] = 238;
assign img[ 2795] = 238;
assign img[ 2796] = 238;
assign img[ 2797] = 238;
assign img[ 2798] = 206;
assign img[ 2799] = 142;
assign img[ 2800] = 136;
assign img[ 2801] = 168;
assign img[ 2802] = 170;
assign img[ 2803] = 238;
assign img[ 2804] = 238;
assign img[ 2805] = 222;
assign img[ 2806] = 253;
assign img[ 2807] = 255;
assign img[ 2808] = 238;
assign img[ 2809] = 254;
assign img[ 2810] = 238;
assign img[ 2811] = 255;
assign img[ 2812] = 238;
assign img[ 2813] = 238;
assign img[ 2814] = 206;
assign img[ 2815] = 238;
assign img[ 2816] = 0;
assign img[ 2817] = 204;
assign img[ 2818] = 236;
assign img[ 2819] = 238;
assign img[ 2820] = 238;
assign img[ 2821] = 238;
assign img[ 2822] = 191;
assign img[ 2823] = 255;
assign img[ 2824] = 255;
assign img[ 2825] = 255;
assign img[ 2826] = 255;
assign img[ 2827] = 239;
assign img[ 2828] = 204;
assign img[ 2829] = 255;
assign img[ 2830] = 255;
assign img[ 2831] = 239;
assign img[ 2832] = 238;
assign img[ 2833] = 238;
assign img[ 2834] = 238;
assign img[ 2835] = 238;
assign img[ 2836] = 238;
assign img[ 2837] = 204;
assign img[ 2838] = 252;
assign img[ 2839] = 255;
assign img[ 2840] = 238;
assign img[ 2841] = 238;
assign img[ 2842] = 238;
assign img[ 2843] = 238;
assign img[ 2844] = 238;
assign img[ 2845] = 255;
assign img[ 2846] = 255;
assign img[ 2847] = 191;
assign img[ 2848] = 251;
assign img[ 2849] = 255;
assign img[ 2850] = 255;
assign img[ 2851] = 255;
assign img[ 2852] = 239;
assign img[ 2853] = 238;
assign img[ 2854] = 238;
assign img[ 2855] = 238;
assign img[ 2856] = 138;
assign img[ 2857] = 238;
assign img[ 2858] = 238;
assign img[ 2859] = 255;
assign img[ 2860] = 238;
assign img[ 2861] = 239;
assign img[ 2862] = 238;
assign img[ 2863] = 238;
assign img[ 2864] = 254;
assign img[ 2865] = 255;
assign img[ 2866] = 255;
assign img[ 2867] = 238;
assign img[ 2868] = 238;
assign img[ 2869] = 238;
assign img[ 2870] = 223;
assign img[ 2871] = 254;
assign img[ 2872] = 255;
assign img[ 2873] = 255;
assign img[ 2874] = 255;
assign img[ 2875] = 255;
assign img[ 2876] = 255;
assign img[ 2877] = 255;
assign img[ 2878] = 255;
assign img[ 2879] = 255;
assign img[ 2880] = 255;
assign img[ 2881] = 239;
assign img[ 2882] = 254;
assign img[ 2883] = 255;
assign img[ 2884] = 255;
assign img[ 2885] = 255;
assign img[ 2886] = 238;
assign img[ 2887] = 238;
assign img[ 2888] = 238;
assign img[ 2889] = 207;
assign img[ 2890] = 238;
assign img[ 2891] = 255;
assign img[ 2892] = 255;
assign img[ 2893] = 239;
assign img[ 2894] = 238;
assign img[ 2895] = 255;
assign img[ 2896] = 255;
assign img[ 2897] = 255;
assign img[ 2898] = 255;
assign img[ 2899] = 255;
assign img[ 2900] = 255;
assign img[ 2901] = 223;
assign img[ 2902] = 253;
assign img[ 2903] = 207;
assign img[ 2904] = 252;
assign img[ 2905] = 239;
assign img[ 2906] = 238;
assign img[ 2907] = 238;
assign img[ 2908] = 255;
assign img[ 2909] = 255;
assign img[ 2910] = 255;
assign img[ 2911] = 255;
assign img[ 2912] = 221;
assign img[ 2913] = 221;
assign img[ 2914] = 253;
assign img[ 2915] = 255;
assign img[ 2916] = 255;
assign img[ 2917] = 223;
assign img[ 2918] = 221;
assign img[ 2919] = 255;
assign img[ 2920] = 239;
assign img[ 2921] = 238;
assign img[ 2922] = 206;
assign img[ 2923] = 220;
assign img[ 2924] = 221;
assign img[ 2925] = 253;
assign img[ 2926] = 255;
assign img[ 2927] = 239;
assign img[ 2928] = 220;
assign img[ 2929] = 236;
assign img[ 2930] = 204;
assign img[ 2931] = 238;
assign img[ 2932] = 206;
assign img[ 2933] = 238;
assign img[ 2934] = 238;
assign img[ 2935] = 238;
assign img[ 2936] = 255;
assign img[ 2937] = 191;
assign img[ 2938] = 255;
assign img[ 2939] = 239;
assign img[ 2940] = 220;
assign img[ 2941] = 255;
assign img[ 2942] = 255;
assign img[ 2943] = 255;
assign img[ 2944] = 96;
assign img[ 2945] = 255;
assign img[ 2946] = 255;
assign img[ 2947] = 255;
assign img[ 2948] = 255;
assign img[ 2949] = 255;
assign img[ 2950] = 255;
assign img[ 2951] = 255;
assign img[ 2952] = 255;
assign img[ 2953] = 255;
assign img[ 2954] = 255;
assign img[ 2955] = 239;
assign img[ 2956] = 138;
assign img[ 2957] = 238;
assign img[ 2958] = 238;
assign img[ 2959] = 206;
assign img[ 2960] = 204;
assign img[ 2961] = 238;
assign img[ 2962] = 206;
assign img[ 2963] = 221;
assign img[ 2964] = 221;
assign img[ 2965] = 253;
assign img[ 2966] = 239;
assign img[ 2967] = 238;
assign img[ 2968] = 238;
assign img[ 2969] = 238;
assign img[ 2970] = 170;
assign img[ 2971] = 238;
assign img[ 2972] = 238;
assign img[ 2973] = 255;
assign img[ 2974] = 255;
assign img[ 2975] = 255;
assign img[ 2976] = 187;
assign img[ 2977] = 255;
assign img[ 2978] = 255;
assign img[ 2979] = 255;
assign img[ 2980] = 255;
assign img[ 2981] = 255;
assign img[ 2982] = 255;
assign img[ 2983] = 255;
assign img[ 2984] = 255;
assign img[ 2985] = 255;
assign img[ 2986] = 255;
assign img[ 2987] = 255;
assign img[ 2988] = 223;
assign img[ 2989] = 221;
assign img[ 2990] = 253;
assign img[ 2991] = 255;
assign img[ 2992] = 238;
assign img[ 2993] = 254;
assign img[ 2994] = 238;
assign img[ 2995] = 255;
assign img[ 2996] = 238;
assign img[ 2997] = 255;
assign img[ 2998] = 238;
assign img[ 2999] = 239;
assign img[ 3000] = 238;
assign img[ 3001] = 254;
assign img[ 3002] = 221;
assign img[ 3003] = 221;
assign img[ 3004] = 255;
assign img[ 3005] = 255;
assign img[ 3006] = 255;
assign img[ 3007] = 255;
assign img[ 3008] = 255;
assign img[ 3009] = 255;
assign img[ 3010] = 239;
assign img[ 3011] = 238;
assign img[ 3012] = 238;
assign img[ 3013] = 238;
assign img[ 3014] = 206;
assign img[ 3015] = 204;
assign img[ 3016] = 204;
assign img[ 3017] = 238;
assign img[ 3018] = 238;
assign img[ 3019] = 254;
assign img[ 3020] = 255;
assign img[ 3021] = 255;
assign img[ 3022] = 255;
assign img[ 3023] = 255;
assign img[ 3024] = 239;
assign img[ 3025] = 238;
assign img[ 3026] = 222;
assign img[ 3027] = 221;
assign img[ 3028] = 253;
assign img[ 3029] = 239;
assign img[ 3030] = 238;
assign img[ 3031] = 238;
assign img[ 3032] = 174;
assign img[ 3033] = 238;
assign img[ 3034] = 238;
assign img[ 3035] = 238;
assign img[ 3036] = 255;
assign img[ 3037] = 255;
assign img[ 3038] = 255;
assign img[ 3039] = 207;
assign img[ 3040] = 236;
assign img[ 3041] = 238;
assign img[ 3042] = 254;
assign img[ 3043] = 255;
assign img[ 3044] = 255;
assign img[ 3045] = 255;
assign img[ 3046] = 191;
assign img[ 3047] = 255;
assign img[ 3048] = 255;
assign img[ 3049] = 255;
assign img[ 3050] = 238;
assign img[ 3051] = 206;
assign img[ 3052] = 204;
assign img[ 3053] = 223;
assign img[ 3054] = 255;
assign img[ 3055] = 239;
assign img[ 3056] = 238;
assign img[ 3057] = 238;
assign img[ 3058] = 254;
assign img[ 3059] = 239;
assign img[ 3060] = 239;
assign img[ 3061] = 238;
assign img[ 3062] = 238;
assign img[ 3063] = 254;
assign img[ 3064] = 254;
assign img[ 3065] = 255;
assign img[ 3066] = 255;
assign img[ 3067] = 255;
assign img[ 3068] = 205;
assign img[ 3069] = 255;
assign img[ 3070] = 255;
assign img[ 3071] = 255;
assign img[ 3072] = 64;
assign img[ 3073] = 204;
assign img[ 3074] = 236;
assign img[ 3075] = 255;
assign img[ 3076] = 255;
assign img[ 3077] = 223;
assign img[ 3078] = 221;
assign img[ 3079] = 255;
assign img[ 3080] = 255;
assign img[ 3081] = 255;
assign img[ 3082] = 238;
assign img[ 3083] = 238;
assign img[ 3084] = 238;
assign img[ 3085] = 238;
assign img[ 3086] = 238;
assign img[ 3087] = 255;
assign img[ 3088] = 206;
assign img[ 3089] = 220;
assign img[ 3090] = 253;
assign img[ 3091] = 174;
assign img[ 3092] = 170;
assign img[ 3093] = 238;
assign img[ 3094] = 238;
assign img[ 3095] = 254;
assign img[ 3096] = 255;
assign img[ 3097] = 191;
assign img[ 3098] = 255;
assign img[ 3099] = 255;
assign img[ 3100] = 255;
assign img[ 3101] = 255;
assign img[ 3102] = 255;
assign img[ 3103] = 255;
assign img[ 3104] = 255;
assign img[ 3105] = 255;
assign img[ 3106] = 255;
assign img[ 3107] = 255;
assign img[ 3108] = 255;
assign img[ 3109] = 255;
assign img[ 3110] = 255;
assign img[ 3111] = 255;
assign img[ 3112] = 255;
assign img[ 3113] = 255;
assign img[ 3114] = 255;
assign img[ 3115] = 255;
assign img[ 3116] = 238;
assign img[ 3117] = 255;
assign img[ 3118] = 238;
assign img[ 3119] = 238;
assign img[ 3120] = 238;
assign img[ 3121] = 239;
assign img[ 3122] = 238;
assign img[ 3123] = 238;
assign img[ 3124] = 238;
assign img[ 3125] = 254;
assign img[ 3126] = 255;
assign img[ 3127] = 238;
assign img[ 3128] = 238;
assign img[ 3129] = 255;
assign img[ 3130] = 239;
assign img[ 3131] = 255;
assign img[ 3132] = 255;
assign img[ 3133] = 255;
assign img[ 3134] = 238;
assign img[ 3135] = 254;
assign img[ 3136] = 255;
assign img[ 3137] = 255;
assign img[ 3138] = 238;
assign img[ 3139] = 238;
assign img[ 3140] = 255;
assign img[ 3141] = 255;
assign img[ 3142] = 255;
assign img[ 3143] = 255;
assign img[ 3144] = 255;
assign img[ 3145] = 255;
assign img[ 3146] = 255;
assign img[ 3147] = 255;
assign img[ 3148] = 238;
assign img[ 3149] = 238;
assign img[ 3150] = 238;
assign img[ 3151] = 238;
assign img[ 3152] = 238;
assign img[ 3153] = 238;
assign img[ 3154] = 238;
assign img[ 3155] = 254;
assign img[ 3156] = 239;
assign img[ 3157] = 238;
assign img[ 3158] = 238;
assign img[ 3159] = 238;
assign img[ 3160] = 222;
assign img[ 3161] = 221;
assign img[ 3162] = 253;
assign img[ 3163] = 255;
assign img[ 3164] = 255;
assign img[ 3165] = 255;
assign img[ 3166] = 255;
assign img[ 3167] = 239;
assign img[ 3168] = 238;
assign img[ 3169] = 223;
assign img[ 3170] = 253;
assign img[ 3171] = 223;
assign img[ 3172] = 253;
assign img[ 3173] = 255;
assign img[ 3174] = 255;
assign img[ 3175] = 255;
assign img[ 3176] = 255;
assign img[ 3177] = 239;
assign img[ 3178] = 238;
assign img[ 3179] = 238;
assign img[ 3180] = 238;
assign img[ 3181] = 238;
assign img[ 3182] = 238;
assign img[ 3183] = 255;
assign img[ 3184] = 204;
assign img[ 3185] = 238;
assign img[ 3186] = 238;
assign img[ 3187] = 238;
assign img[ 3188] = 206;
assign img[ 3189] = 220;
assign img[ 3190] = 205;
assign img[ 3191] = 236;
assign img[ 3192] = 238;
assign img[ 3193] = 238;
assign img[ 3194] = 138;
assign img[ 3195] = 136;
assign img[ 3196] = 200;
assign img[ 3197] = 238;
assign img[ 3198] = 238;
assign img[ 3199] = 238;
assign img[ 3200] = 96;
assign img[ 3201] = 255;
assign img[ 3202] = 255;
assign img[ 3203] = 255;
assign img[ 3204] = 223;
assign img[ 3205] = 205;
assign img[ 3206] = 252;
assign img[ 3207] = 255;
assign img[ 3208] = 255;
assign img[ 3209] = 255;
assign img[ 3210] = 255;
assign img[ 3211] = 255;
assign img[ 3212] = 238;
assign img[ 3213] = 238;
assign img[ 3214] = 238;
assign img[ 3215] = 207;
assign img[ 3216] = 204;
assign img[ 3217] = 236;
assign img[ 3218] = 238;
assign img[ 3219] = 238;
assign img[ 3220] = 254;
assign img[ 3221] = 255;
assign img[ 3222] = 255;
assign img[ 3223] = 255;
assign img[ 3224] = 255;
assign img[ 3225] = 207;
assign img[ 3226] = 204;
assign img[ 3227] = 238;
assign img[ 3228] = 238;
assign img[ 3229] = 238;
assign img[ 3230] = 254;
assign img[ 3231] = 255;
assign img[ 3232] = 170;
assign img[ 3233] = 239;
assign img[ 3234] = 254;
assign img[ 3235] = 255;
assign img[ 3236] = 255;
assign img[ 3237] = 255;
assign img[ 3238] = 255;
assign img[ 3239] = 207;
assign img[ 3240] = 236;
assign img[ 3241] = 238;
assign img[ 3242] = 238;
assign img[ 3243] = 238;
assign img[ 3244] = 220;
assign img[ 3245] = 221;
assign img[ 3246] = 253;
assign img[ 3247] = 207;
assign img[ 3248] = 236;
assign img[ 3249] = 238;
assign img[ 3250] = 238;
assign img[ 3251] = 238;
assign img[ 3252] = 254;
assign img[ 3253] = 255;
assign img[ 3254] = 255;
assign img[ 3255] = 255;
assign img[ 3256] = 255;
assign img[ 3257] = 255;
assign img[ 3258] = 255;
assign img[ 3259] = 255;
assign img[ 3260] = 255;
assign img[ 3261] = 239;
assign img[ 3262] = 204;
assign img[ 3263] = 238;
assign img[ 3264] = 238;
assign img[ 3265] = 238;
assign img[ 3266] = 254;
assign img[ 3267] = 254;
assign img[ 3268] = 238;
assign img[ 3269] = 255;
assign img[ 3270] = 204;
assign img[ 3271] = 252;
assign img[ 3272] = 255;
assign img[ 3273] = 255;
assign img[ 3274] = 238;
assign img[ 3275] = 254;
assign img[ 3276] = 255;
assign img[ 3277] = 255;
assign img[ 3278] = 255;
assign img[ 3279] = 255;
assign img[ 3280] = 223;
assign img[ 3281] = 255;
assign img[ 3282] = 255;
assign img[ 3283] = 255;
assign img[ 3284] = 223;
assign img[ 3285] = 221;
assign img[ 3286] = 253;
assign img[ 3287] = 255;
assign img[ 3288] = 191;
assign img[ 3289] = 255;
assign img[ 3290] = 223;
assign img[ 3291] = 255;
assign img[ 3292] = 255;
assign img[ 3293] = 255;
assign img[ 3294] = 255;
assign img[ 3295] = 223;
assign img[ 3296] = 255;
assign img[ 3297] = 239;
assign img[ 3298] = 238;
assign img[ 3299] = 255;
assign img[ 3300] = 255;
assign img[ 3301] = 255;
assign img[ 3302] = 223;
assign img[ 3303] = 255;
assign img[ 3304] = 255;
assign img[ 3305] = 255;
assign img[ 3306] = 238;
assign img[ 3307] = 238;
assign img[ 3308] = 238;
assign img[ 3309] = 238;
assign img[ 3310] = 238;
assign img[ 3311] = 238;
assign img[ 3312] = 238;
assign img[ 3313] = 238;
assign img[ 3314] = 238;
assign img[ 3315] = 206;
assign img[ 3316] = 204;
assign img[ 3317] = 236;
assign img[ 3318] = 238;
assign img[ 3319] = 238;
assign img[ 3320] = 238;
assign img[ 3321] = 206;
assign img[ 3322] = 204;
assign img[ 3323] = 204;
assign img[ 3324] = 236;
assign img[ 3325] = 238;
assign img[ 3326] = 238;
assign img[ 3327] = 238;
assign img[ 3328] = 96;
assign img[ 3329] = 207;
assign img[ 3330] = 236;
assign img[ 3331] = 206;
assign img[ 3332] = 236;
assign img[ 3333] = 254;
assign img[ 3334] = 191;
assign img[ 3335] = 255;
assign img[ 3336] = 255;
assign img[ 3337] = 239;
assign img[ 3338] = 238;
assign img[ 3339] = 255;
assign img[ 3340] = 255;
assign img[ 3341] = 255;
assign img[ 3342] = 255;
assign img[ 3343] = 255;
assign img[ 3344] = 187;
assign img[ 3345] = 251;
assign img[ 3346] = 255;
assign img[ 3347] = 255;
assign img[ 3348] = 153;
assign img[ 3349] = 187;
assign img[ 3350] = 255;
assign img[ 3351] = 239;
assign img[ 3352] = 238;
assign img[ 3353] = 255;
assign img[ 3354] = 221;
assign img[ 3355] = 253;
assign img[ 3356] = 255;
assign img[ 3357] = 255;
assign img[ 3358] = 239;
assign img[ 3359] = 238;
assign img[ 3360] = 238;
assign img[ 3361] = 255;
assign img[ 3362] = 175;
assign img[ 3363] = 238;
assign img[ 3364] = 238;
assign img[ 3365] = 238;
assign img[ 3366] = 238;
assign img[ 3367] = 255;
assign img[ 3368] = 255;
assign img[ 3369] = 255;
assign img[ 3370] = 239;
assign img[ 3371] = 238;
assign img[ 3372] = 238;
assign img[ 3373] = 238;
assign img[ 3374] = 238;
assign img[ 3375] = 223;
assign img[ 3376] = 253;
assign img[ 3377] = 255;
assign img[ 3378] = 255;
assign img[ 3379] = 255;
assign img[ 3380] = 255;
assign img[ 3381] = 255;
assign img[ 3382] = 255;
assign img[ 3383] = 255;
assign img[ 3384] = 221;
assign img[ 3385] = 255;
assign img[ 3386] = 255;
assign img[ 3387] = 255;
assign img[ 3388] = 255;
assign img[ 3389] = 191;
assign img[ 3390] = 255;
assign img[ 3391] = 255;
assign img[ 3392] = 255;
assign img[ 3393] = 255;
assign img[ 3394] = 255;
assign img[ 3395] = 255;
assign img[ 3396] = 255;
assign img[ 3397] = 255;
assign img[ 3398] = 255;
assign img[ 3399] = 255;
assign img[ 3400] = 238;
assign img[ 3401] = 238;
assign img[ 3402] = 255;
assign img[ 3403] = 255;
assign img[ 3404] = 205;
assign img[ 3405] = 204;
assign img[ 3406] = 238;
assign img[ 3407] = 255;
assign img[ 3408] = 255;
assign img[ 3409] = 255;
assign img[ 3410] = 223;
assign img[ 3411] = 255;
assign img[ 3412] = 255;
assign img[ 3413] = 223;
assign img[ 3414] = 238;
assign img[ 3415] = 238;
assign img[ 3416] = 174;
assign img[ 3417] = 254;
assign img[ 3418] = 238;
assign img[ 3419] = 238;
assign img[ 3420] = 238;
assign img[ 3421] = 175;
assign img[ 3422] = 255;
assign img[ 3423] = 255;
assign img[ 3424] = 255;
assign img[ 3425] = 255;
assign img[ 3426] = 238;
assign img[ 3427] = 238;
assign img[ 3428] = 238;
assign img[ 3429] = 255;
assign img[ 3430] = 221;
assign img[ 3431] = 253;
assign img[ 3432] = 255;
assign img[ 3433] = 255;
assign img[ 3434] = 255;
assign img[ 3435] = 255;
assign img[ 3436] = 238;
assign img[ 3437] = 238;
assign img[ 3438] = 254;
assign img[ 3439] = 239;
assign img[ 3440] = 254;
assign img[ 3441] = 255;
assign img[ 3442] = 255;
assign img[ 3443] = 255;
assign img[ 3444] = 255;
assign img[ 3445] = 239;
assign img[ 3446] = 238;
assign img[ 3447] = 255;
assign img[ 3448] = 255;
assign img[ 3449] = 191;
assign img[ 3450] = 185;
assign img[ 3451] = 171;
assign img[ 3452] = 250;
assign img[ 3453] = 255;
assign img[ 3454] = 239;
assign img[ 3455] = 238;
assign img[ 3456] = 80;
assign img[ 3457] = 101;
assign img[ 3458] = 118;
assign img[ 3459] = 207;
assign img[ 3460] = 204;
assign img[ 3461] = 204;
assign img[ 3462] = 204;
assign img[ 3463] = 236;
assign img[ 3464] = 238;
assign img[ 3465] = 238;
assign img[ 3466] = 238;
assign img[ 3467] = 255;
assign img[ 3468] = 255;
assign img[ 3469] = 255;
assign img[ 3470] = 255;
assign img[ 3471] = 223;
assign img[ 3472] = 221;
assign img[ 3473] = 221;
assign img[ 3474] = 253;
assign img[ 3475] = 191;
assign img[ 3476] = 187;
assign img[ 3477] = 255;
assign img[ 3478] = 255;
assign img[ 3479] = 255;
assign img[ 3480] = 255;
assign img[ 3481] = 255;
assign img[ 3482] = 239;
assign img[ 3483] = 238;
assign img[ 3484] = 238;
assign img[ 3485] = 238;
assign img[ 3486] = 254;
assign img[ 3487] = 255;
assign img[ 3488] = 255;
assign img[ 3489] = 255;
assign img[ 3490] = 255;
assign img[ 3491] = 255;
assign img[ 3492] = 255;
assign img[ 3493] = 255;
assign img[ 3494] = 239;
assign img[ 3495] = 239;
assign img[ 3496] = 238;
assign img[ 3497] = 238;
assign img[ 3498] = 254;
assign img[ 3499] = 255;
assign img[ 3500] = 238;
assign img[ 3501] = 238;
assign img[ 3502] = 238;
assign img[ 3503] = 238;
assign img[ 3504] = 254;
assign img[ 3505] = 255;
assign img[ 3506] = 255;
assign img[ 3507] = 255;
assign img[ 3508] = 239;
assign img[ 3509] = 255;
assign img[ 3510] = 255;
assign img[ 3511] = 191;
assign img[ 3512] = 187;
assign img[ 3513] = 255;
assign img[ 3514] = 255;
assign img[ 3515] = 255;
assign img[ 3516] = 255;
assign img[ 3517] = 239;
assign img[ 3518] = 238;
assign img[ 3519] = 255;
assign img[ 3520] = 255;
assign img[ 3521] = 255;
assign img[ 3522] = 255;
assign img[ 3523] = 255;
assign img[ 3524] = 255;
assign img[ 3525] = 255;
assign img[ 3526] = 255;
assign img[ 3527] = 255;
assign img[ 3528] = 221;
assign img[ 3529] = 255;
assign img[ 3530] = 255;
assign img[ 3531] = 239;
assign img[ 3532] = 238;
assign img[ 3533] = 238;
assign img[ 3534] = 238;
assign img[ 3535] = 255;
assign img[ 3536] = 239;
assign img[ 3537] = 238;
assign img[ 3538] = 206;
assign img[ 3539] = 238;
assign img[ 3540] = 238;
assign img[ 3541] = 238;
assign img[ 3542] = 238;
assign img[ 3543] = 238;
assign img[ 3544] = 206;
assign img[ 3545] = 204;
assign img[ 3546] = 236;
assign img[ 3547] = 238;
assign img[ 3548] = 238;
assign img[ 3549] = 238;
assign img[ 3550] = 238;
assign img[ 3551] = 174;
assign img[ 3552] = 238;
assign img[ 3553] = 238;
assign img[ 3554] = 238;
assign img[ 3555] = 239;
assign img[ 3556] = 254;
assign img[ 3557] = 223;
assign img[ 3558] = 255;
assign img[ 3559] = 255;
assign img[ 3560] = 255;
assign img[ 3561] = 255;
assign img[ 3562] = 255;
assign img[ 3563] = 255;
assign img[ 3564] = 191;
assign img[ 3565] = 255;
assign img[ 3566] = 255;
assign img[ 3567] = 255;
assign img[ 3568] = 255;
assign img[ 3569] = 255;
assign img[ 3570] = 223;
assign img[ 3571] = 221;
assign img[ 3572] = 253;
assign img[ 3573] = 255;
assign img[ 3574] = 255;
assign img[ 3575] = 255;
assign img[ 3576] = 255;
assign img[ 3577] = 255;
assign img[ 3578] = 187;
assign img[ 3579] = 153;
assign img[ 3580] = 153;
assign img[ 3581] = 253;
assign img[ 3582] = 255;
assign img[ 3583] = 255;
assign img[ 3584] = 32;
assign img[ 3585] = 138;
assign img[ 3586] = 232;
assign img[ 3587] = 238;
assign img[ 3588] = 254;
assign img[ 3589] = 255;
assign img[ 3590] = 255;
assign img[ 3591] = 255;
assign img[ 3592] = 238;
assign img[ 3593] = 238;
assign img[ 3594] = 238;
assign img[ 3595] = 238;
assign img[ 3596] = 206;
assign img[ 3597] = 220;
assign img[ 3598] = 205;
assign img[ 3599] = 204;
assign img[ 3600] = 236;
assign img[ 3601] = 238;
assign img[ 3602] = 238;
assign img[ 3603] = 255;
assign img[ 3604] = 238;
assign img[ 3605] = 254;
assign img[ 3606] = 239;
assign img[ 3607] = 238;
assign img[ 3608] = 238;
assign img[ 3609] = 207;
assign img[ 3610] = 204;
assign img[ 3611] = 220;
assign img[ 3612] = 253;
assign img[ 3613] = 255;
assign img[ 3614] = 223;
assign img[ 3615] = 221;
assign img[ 3616] = 204;
assign img[ 3617] = 236;
assign img[ 3618] = 238;
assign img[ 3619] = 255;
assign img[ 3620] = 255;
assign img[ 3621] = 255;
assign img[ 3622] = 255;
assign img[ 3623] = 255;
assign img[ 3624] = 255;
assign img[ 3625] = 255;
assign img[ 3626] = 238;
assign img[ 3627] = 238;
assign img[ 3628] = 238;
assign img[ 3629] = 206;
assign img[ 3630] = 238;
assign img[ 3631] = 255;
assign img[ 3632] = 255;
assign img[ 3633] = 255;
assign img[ 3634] = 255;
assign img[ 3635] = 255;
assign img[ 3636] = 239;
assign img[ 3637] = 255;
assign img[ 3638] = 255;
assign img[ 3639] = 255;
assign img[ 3640] = 255;
assign img[ 3641] = 255;
assign img[ 3642] = 255;
assign img[ 3643] = 255;
assign img[ 3644] = 255;
assign img[ 3645] = 255;
assign img[ 3646] = 255;
assign img[ 3647] = 255;
assign img[ 3648] = 255;
assign img[ 3649] = 255;
assign img[ 3650] = 223;
assign img[ 3651] = 255;
assign img[ 3652] = 255;
assign img[ 3653] = 255;
assign img[ 3654] = 239;
assign img[ 3655] = 238;
assign img[ 3656] = 238;
assign img[ 3657] = 238;
assign img[ 3658] = 254;
assign img[ 3659] = 223;
assign img[ 3660] = 204;
assign img[ 3661] = 238;
assign img[ 3662] = 238;
assign img[ 3663] = 255;
assign img[ 3664] = 239;
assign img[ 3665] = 238;
assign img[ 3666] = 238;
assign img[ 3667] = 238;
assign img[ 3668] = 254;
assign img[ 3669] = 255;
assign img[ 3670] = 238;
assign img[ 3671] = 238;
assign img[ 3672] = 254;
assign img[ 3673] = 255;
assign img[ 3674] = 255;
assign img[ 3675] = 255;
assign img[ 3676] = 255;
assign img[ 3677] = 255;
assign img[ 3678] = 255;
assign img[ 3679] = 223;
assign img[ 3680] = 204;
assign img[ 3681] = 204;
assign img[ 3682] = 252;
assign img[ 3683] = 255;
assign img[ 3684] = 223;
assign img[ 3685] = 221;
assign img[ 3686] = 136;
assign img[ 3687] = 136;
assign img[ 3688] = 236;
assign img[ 3689] = 238;
assign img[ 3690] = 254;
assign img[ 3691] = 255;
assign img[ 3692] = 238;
assign img[ 3693] = 238;
assign img[ 3694] = 238;
assign img[ 3695] = 238;
assign img[ 3696] = 238;
assign img[ 3697] = 206;
assign img[ 3698] = 204;
assign img[ 3699] = 204;
assign img[ 3700] = 253;
assign img[ 3701] = 238;
assign img[ 3702] = 238;
assign img[ 3703] = 254;
assign img[ 3704] = 238;
assign img[ 3705] = 238;
assign img[ 3706] = 238;
assign img[ 3707] = 238;
assign img[ 3708] = 238;
assign img[ 3709] = 238;
assign img[ 3710] = 222;
assign img[ 3711] = 221;
assign img[ 3712] = 96;
assign img[ 3713] = 206;
assign img[ 3714] = 204;
assign img[ 3715] = 204;
assign img[ 3716] = 204;
assign img[ 3717] = 238;
assign img[ 3718] = 254;
assign img[ 3719] = 255;
assign img[ 3720] = 238;
assign img[ 3721] = 238;
assign img[ 3722] = 190;
assign img[ 3723] = 187;
assign img[ 3724] = 251;
assign img[ 3725] = 255;
assign img[ 3726] = 255;
assign img[ 3727] = 191;
assign img[ 3728] = 251;
assign img[ 3729] = 223;
assign img[ 3730] = 253;
assign img[ 3731] = 191;
assign img[ 3732] = 187;
assign img[ 3733] = 255;
assign img[ 3734] = 223;
assign img[ 3735] = 255;
assign img[ 3736] = 255;
assign img[ 3737] = 255;
assign img[ 3738] = 255;
assign img[ 3739] = 255;
assign img[ 3740] = 255;
assign img[ 3741] = 255;
assign img[ 3742] = 255;
assign img[ 3743] = 191;
assign img[ 3744] = 251;
assign img[ 3745] = 255;
assign img[ 3746] = 255;
assign img[ 3747] = 255;
assign img[ 3748] = 255;
assign img[ 3749] = 255;
assign img[ 3750] = 255;
assign img[ 3751] = 255;
assign img[ 3752] = 255;
assign img[ 3753] = 255;
assign img[ 3754] = 239;
assign img[ 3755] = 238;
assign img[ 3756] = 254;
assign img[ 3757] = 255;
assign img[ 3758] = 255;
assign img[ 3759] = 223;
assign img[ 3760] = 255;
assign img[ 3761] = 255;
assign img[ 3762] = 255;
assign img[ 3763] = 239;
assign img[ 3764] = 238;
assign img[ 3765] = 238;
assign img[ 3766] = 191;
assign img[ 3767] = 255;
assign img[ 3768] = 255;
assign img[ 3769] = 255;
assign img[ 3770] = 223;
assign img[ 3771] = 255;
assign img[ 3772] = 254;
assign img[ 3773] = 223;
assign img[ 3774] = 254;
assign img[ 3775] = 254;
assign img[ 3776] = 238;
assign img[ 3777] = 255;
assign img[ 3778] = 254;
assign img[ 3779] = 255;
assign img[ 3780] = 255;
assign img[ 3781] = 255;
assign img[ 3782] = 238;
assign img[ 3783] = 238;
assign img[ 3784] = 238;
assign img[ 3785] = 254;
assign img[ 3786] = 238;
assign img[ 3787] = 238;
assign img[ 3788] = 238;
assign img[ 3789] = 238;
assign img[ 3790] = 238;
assign img[ 3791] = 255;
assign img[ 3792] = 223;
assign img[ 3793] = 255;
assign img[ 3794] = 191;
assign img[ 3795] = 255;
assign img[ 3796] = 239;
assign img[ 3797] = 255;
assign img[ 3798] = 255;
assign img[ 3799] = 255;
assign img[ 3800] = 223;
assign img[ 3801] = 221;
assign img[ 3802] = 221;
assign img[ 3803] = 221;
assign img[ 3804] = 253;
assign img[ 3805] = 255;
assign img[ 3806] = 255;
assign img[ 3807] = 255;
assign img[ 3808] = 221;
assign img[ 3809] = 221;
assign img[ 3810] = 253;
assign img[ 3811] = 255;
assign img[ 3812] = 255;
assign img[ 3813] = 239;
assign img[ 3814] = 238;
assign img[ 3815] = 238;
assign img[ 3816] = 254;
assign img[ 3817] = 239;
assign img[ 3818] = 238;
assign img[ 3819] = 238;
assign img[ 3820] = 254;
assign img[ 3821] = 255;
assign img[ 3822] = 255;
assign img[ 3823] = 223;
assign img[ 3824] = 172;
assign img[ 3825] = 187;
assign img[ 3826] = 251;
assign img[ 3827] = 255;
assign img[ 3828] = 221;
assign img[ 3829] = 191;
assign img[ 3830] = 251;
assign img[ 3831] = 255;
assign img[ 3832] = 239;
assign img[ 3833] = 238;
assign img[ 3834] = 238;
assign img[ 3835] = 238;
assign img[ 3836] = 254;
assign img[ 3837] = 255;
assign img[ 3838] = 223;
assign img[ 3839] = 255;
assign img[ 3840] = 96;
assign img[ 3841] = 255;
assign img[ 3842] = 255;
assign img[ 3843] = 255;
assign img[ 3844] = 253;
assign img[ 3845] = 253;
assign img[ 3846] = 253;
assign img[ 3847] = 255;
assign img[ 3848] = 255;
assign img[ 3849] = 255;
assign img[ 3850] = 255;
assign img[ 3851] = 255;
assign img[ 3852] = 221;
assign img[ 3853] = 255;
assign img[ 3854] = 239;
assign img[ 3855] = 238;
assign img[ 3856] = 238;
assign img[ 3857] = 238;
assign img[ 3858] = 254;
assign img[ 3859] = 255;
assign img[ 3860] = 255;
assign img[ 3861] = 255;
assign img[ 3862] = 223;
assign img[ 3863] = 255;
assign img[ 3864] = 255;
assign img[ 3865] = 255;
assign img[ 3866] = 155;
assign img[ 3867] = 255;
assign img[ 3868] = 255;
assign img[ 3869] = 255;
assign img[ 3870] = 255;
assign img[ 3871] = 191;
assign img[ 3872] = 138;
assign img[ 3873] = 255;
assign img[ 3874] = 255;
assign img[ 3875] = 255;
assign img[ 3876] = 255;
assign img[ 3877] = 255;
assign img[ 3878] = 255;
assign img[ 3879] = 255;
assign img[ 3880] = 255;
assign img[ 3881] = 255;
assign img[ 3882] = 255;
assign img[ 3883] = 159;
assign img[ 3884] = 153;
assign img[ 3885] = 155;
assign img[ 3886] = 251;
assign img[ 3887] = 255;
assign img[ 3888] = 255;
assign img[ 3889] = 255;
assign img[ 3890] = 255;
assign img[ 3891] = 255;
assign img[ 3892] = 255;
assign img[ 3893] = 255;
assign img[ 3894] = 255;
assign img[ 3895] = 255;
assign img[ 3896] = 255;
assign img[ 3897] = 255;
assign img[ 3898] = 239;
assign img[ 3899] = 238;
assign img[ 3900] = 238;
assign img[ 3901] = 206;
assign img[ 3902] = 204;
assign img[ 3903] = 255;
assign img[ 3904] = 255;
assign img[ 3905] = 255;
assign img[ 3906] = 223;
assign img[ 3907] = 255;
assign img[ 3908] = 255;
assign img[ 3909] = 239;
assign img[ 3910] = 238;
assign img[ 3911] = 238;
assign img[ 3912] = 238;
assign img[ 3913] = 238;
assign img[ 3914] = 254;
assign img[ 3915] = 255;
assign img[ 3916] = 191;
assign img[ 3917] = 255;
assign img[ 3918] = 255;
assign img[ 3919] = 255;
assign img[ 3920] = 255;
assign img[ 3921] = 255;
assign img[ 3922] = 223;
assign img[ 3923] = 255;
assign img[ 3924] = 159;
assign img[ 3925] = 253;
assign img[ 3926] = 238;
assign img[ 3927] = 238;
assign img[ 3928] = 206;
assign img[ 3929] = 204;
assign img[ 3930] = 204;
assign img[ 3931] = 204;
assign img[ 3932] = 236;
assign img[ 3933] = 238;
assign img[ 3934] = 254;
assign img[ 3935] = 223;
assign img[ 3936] = 205;
assign img[ 3937] = 255;
assign img[ 3938] = 255;
assign img[ 3939] = 255;
assign img[ 3940] = 255;
assign img[ 3941] = 255;
assign img[ 3942] = 255;
assign img[ 3943] = 255;
assign img[ 3944] = 255;
assign img[ 3945] = 255;
assign img[ 3946] = 255;
assign img[ 3947] = 255;
assign img[ 3948] = 255;
assign img[ 3949] = 255;
assign img[ 3950] = 255;
assign img[ 3951] = 255;
assign img[ 3952] = 255;
assign img[ 3953] = 255;
assign img[ 3954] = 238;
assign img[ 3955] = 238;
assign img[ 3956] = 238;
assign img[ 3957] = 238;
assign img[ 3958] = 238;
assign img[ 3959] = 238;
assign img[ 3960] = 238;
assign img[ 3961] = 255;
assign img[ 3962] = 170;
assign img[ 3963] = 254;
assign img[ 3964] = 254;
assign img[ 3965] = 255;
assign img[ 3966] = 255;
assign img[ 3967] = 255;
assign img[ 3968] = 96;
assign img[ 3969] = 255;
assign img[ 3970] = 255;
assign img[ 3971] = 223;
assign img[ 3972] = 221;
assign img[ 3973] = 221;
assign img[ 3974] = 221;
assign img[ 3975] = 253;
assign img[ 3976] = 255;
assign img[ 3977] = 255;
assign img[ 3978] = 255;
assign img[ 3979] = 255;
assign img[ 3980] = 255;
assign img[ 3981] = 255;
assign img[ 3982] = 255;
assign img[ 3983] = 239;
assign img[ 3984] = 238;
assign img[ 3985] = 255;
assign img[ 3986] = 255;
assign img[ 3987] = 255;
assign img[ 3988] = 171;
assign img[ 3989] = 251;
assign img[ 3990] = 255;
assign img[ 3991] = 255;
assign img[ 3992] = 255;
assign img[ 3993] = 255;
assign img[ 3994] = 238;
assign img[ 3995] = 238;
assign img[ 3996] = 238;
assign img[ 3997] = 238;
assign img[ 3998] = 254;
assign img[ 3999] = 223;
assign img[ 4000] = 237;
assign img[ 4001] = 238;
assign img[ 4002] = 238;
assign img[ 4003] = 255;
assign img[ 4004] = 239;
assign img[ 4005] = 238;
assign img[ 4006] = 238;
assign img[ 4007] = 238;
assign img[ 4008] = 238;
assign img[ 4009] = 238;
assign img[ 4010] = 254;
assign img[ 4011] = 255;
assign img[ 4012] = 191;
assign img[ 4013] = 255;
assign img[ 4014] = 254;
assign img[ 4015] = 238;
assign img[ 4016] = 238;
assign img[ 4017] = 238;
assign img[ 4018] = 238;
assign img[ 4019] = 238;
assign img[ 4020] = 238;
assign img[ 4021] = 254;
assign img[ 4022] = 255;
assign img[ 4023] = 238;
assign img[ 4024] = 238;
assign img[ 4025] = 238;
assign img[ 4026] = 254;
assign img[ 4027] = 255;
assign img[ 4028] = 255;
assign img[ 4029] = 255;
assign img[ 4030] = 255;
assign img[ 4031] = 255;
assign img[ 4032] = 255;
assign img[ 4033] = 255;
assign img[ 4034] = 255;
assign img[ 4035] = 255;
assign img[ 4036] = 255;
assign img[ 4037] = 223;
assign img[ 4038] = 221;
assign img[ 4039] = 255;
assign img[ 4040] = 255;
assign img[ 4041] = 239;
assign img[ 4042] = 238;
assign img[ 4043] = 238;
assign img[ 4044] = 238;
assign img[ 4045] = 238;
assign img[ 4046] = 238;
assign img[ 4047] = 254;
assign img[ 4048] = 255;
assign img[ 4049] = 254;
assign img[ 4050] = 223;
assign img[ 4051] = 157;
assign img[ 4052] = 185;
assign img[ 4053] = 187;
assign img[ 4054] = 234;
assign img[ 4055] = 238;
assign img[ 4056] = 223;
assign img[ 4057] = 255;
assign img[ 4058] = 255;
assign img[ 4059] = 255;
assign img[ 4060] = 255;
assign img[ 4061] = 255;
assign img[ 4062] = 255;
assign img[ 4063] = 239;
assign img[ 4064] = 238;
assign img[ 4065] = 255;
assign img[ 4066] = 255;
assign img[ 4067] = 255;
assign img[ 4068] = 255;
assign img[ 4069] = 239;
assign img[ 4070] = 238;
assign img[ 4071] = 238;
assign img[ 4072] = 254;
assign img[ 4073] = 255;
assign img[ 4074] = 204;
assign img[ 4075] = 204;
assign img[ 4076] = 204;
assign img[ 4077] = 236;
assign img[ 4078] = 238;
assign img[ 4079] = 238;
assign img[ 4080] = 206;
assign img[ 4081] = 238;
assign img[ 4082] = 238;
assign img[ 4083] = 238;
assign img[ 4084] = 238;
assign img[ 4085] = 238;
assign img[ 4086] = 238;
assign img[ 4087] = 238;
assign img[ 4088] = 238;
assign img[ 4089] = 238;
assign img[ 4090] = 238;
assign img[ 4091] = 206;
assign img[ 4092] = 204;
assign img[ 4093] = 236;
assign img[ 4094] = 238;
assign img[ 4095] = 238;
assign img[ 4096] = 96;
assign img[ 4097] = 255;
assign img[ 4098] = 255;
assign img[ 4099] = 223;
assign img[ 4100] = 221;
assign img[ 4101] = 253;
assign img[ 4102] = 255;
assign img[ 4103] = 223;
assign img[ 4104] = 236;
assign img[ 4105] = 254;
assign img[ 4106] = 238;
assign img[ 4107] = 206;
assign img[ 4108] = 220;
assign img[ 4109] = 221;
assign img[ 4110] = 221;
assign img[ 4111] = 221;
assign img[ 4112] = 221;
assign img[ 4113] = 221;
assign img[ 4114] = 253;
assign img[ 4115] = 255;
assign img[ 4116] = 238;
assign img[ 4117] = 238;
assign img[ 4118] = 255;
assign img[ 4119] = 255;
assign img[ 4120] = 238;
assign img[ 4121] = 238;
assign img[ 4122] = 206;
assign img[ 4123] = 238;
assign img[ 4124] = 238;
assign img[ 4125] = 238;
assign img[ 4126] = 238;
assign img[ 4127] = 174;
assign img[ 4128] = 170;
assign img[ 4129] = 238;
assign img[ 4130] = 238;
assign img[ 4131] = 255;
assign img[ 4132] = 239;
assign img[ 4133] = 238;
assign img[ 4134] = 238;
assign img[ 4135] = 238;
assign img[ 4136] = 238;
assign img[ 4137] = 238;
assign img[ 4138] = 238;
assign img[ 4139] = 238;
assign img[ 4140] = 254;
assign img[ 4141] = 255;
assign img[ 4142] = 238;
assign img[ 4143] = 206;
assign img[ 4144] = 254;
assign img[ 4145] = 255;
assign img[ 4146] = 255;
assign img[ 4147] = 255;
assign img[ 4148] = 221;
assign img[ 4149] = 253;
assign img[ 4150] = 254;
assign img[ 4151] = 255;
assign img[ 4152] = 255;
assign img[ 4153] = 255;
assign img[ 4154] = 255;
assign img[ 4155] = 255;
assign img[ 4156] = 255;
assign img[ 4157] = 255;
assign img[ 4158] = 255;
assign img[ 4159] = 255;
assign img[ 4160] = 255;
assign img[ 4161] = 255;
assign img[ 4162] = 223;
assign img[ 4163] = 255;
assign img[ 4164] = 255;
assign img[ 4165] = 239;
assign img[ 4166] = 254;
assign img[ 4167] = 223;
assign img[ 4168] = 253;
assign img[ 4169] = 255;
assign img[ 4170] = 255;
assign img[ 4171] = 255;
assign img[ 4172] = 255;
assign img[ 4173] = 255;
assign img[ 4174] = 238;
assign img[ 4175] = 255;
assign img[ 4176] = 223;
assign img[ 4177] = 255;
assign img[ 4178] = 255;
assign img[ 4179] = 255;
assign img[ 4180] = 255;
assign img[ 4181] = 255;
assign img[ 4182] = 238;
assign img[ 4183] = 255;
assign img[ 4184] = 255;
assign img[ 4185] = 255;
assign img[ 4186] = 222;
assign img[ 4187] = 221;
assign img[ 4188] = 253;
assign img[ 4189] = 255;
assign img[ 4190] = 255;
assign img[ 4191] = 255;
assign img[ 4192] = 191;
assign img[ 4193] = 187;
assign img[ 4194] = 251;
assign img[ 4195] = 239;
assign img[ 4196] = 238;
assign img[ 4197] = 255;
assign img[ 4198] = 221;
assign img[ 4199] = 255;
assign img[ 4200] = 255;
assign img[ 4201] = 239;
assign img[ 4202] = 238;
assign img[ 4203] = 238;
assign img[ 4204] = 238;
assign img[ 4205] = 238;
assign img[ 4206] = 254;
assign img[ 4207] = 223;
assign img[ 4208] = 221;
assign img[ 4209] = 253;
assign img[ 4210] = 206;
assign img[ 4211] = 220;
assign img[ 4212] = 204;
assign img[ 4213] = 204;
assign img[ 4214] = 236;
assign img[ 4215] = 238;
assign img[ 4216] = 238;
assign img[ 4217] = 174;
assign img[ 4218] = 238;
assign img[ 4219] = 206;
assign img[ 4220] = 220;
assign img[ 4221] = 253;
assign img[ 4222] = 223;
assign img[ 4223] = 253;
assign img[ 4224] = 96;
assign img[ 4225] = 239;
assign img[ 4226] = 238;
assign img[ 4227] = 238;
assign img[ 4228] = 206;
assign img[ 4229] = 238;
assign img[ 4230] = 238;
assign img[ 4231] = 254;
assign img[ 4232] = 255;
assign img[ 4233] = 255;
assign img[ 4234] = 255;
assign img[ 4235] = 255;
assign img[ 4236] = 221;
assign img[ 4237] = 253;
assign img[ 4238] = 223;
assign img[ 4239] = 189;
assign img[ 4240] = 255;
assign img[ 4241] = 255;
assign img[ 4242] = 239;
assign img[ 4243] = 238;
assign img[ 4244] = 204;
assign img[ 4245] = 238;
assign img[ 4246] = 206;
assign img[ 4247] = 255;
assign img[ 4248] = 255;
assign img[ 4249] = 255;
assign img[ 4250] = 204;
assign img[ 4251] = 236;
assign img[ 4252] = 238;
assign img[ 4253] = 255;
assign img[ 4254] = 255;
assign img[ 4255] = 255;
assign img[ 4256] = 221;
assign img[ 4257] = 253;
assign img[ 4258] = 255;
assign img[ 4259] = 255;
assign img[ 4260] = 255;
assign img[ 4261] = 255;
assign img[ 4262] = 255;
assign img[ 4263] = 223;
assign img[ 4264] = 221;
assign img[ 4265] = 223;
assign img[ 4266] = 236;
assign img[ 4267] = 254;
assign img[ 4268] = 255;
assign img[ 4269] = 255;
assign img[ 4270] = 255;
assign img[ 4271] = 255;
assign img[ 4272] = 255;
assign img[ 4273] = 255;
assign img[ 4274] = 255;
assign img[ 4275] = 255;
assign img[ 4276] = 255;
assign img[ 4277] = 255;
assign img[ 4278] = 255;
assign img[ 4279] = 255;
assign img[ 4280] = 255;
assign img[ 4281] = 255;
assign img[ 4282] = 223;
assign img[ 4283] = 223;
assign img[ 4284] = 255;
assign img[ 4285] = 255;
assign img[ 4286] = 255;
assign img[ 4287] = 255;
assign img[ 4288] = 255;
assign img[ 4289] = 255;
assign img[ 4290] = 223;
assign img[ 4291] = 255;
assign img[ 4292] = 223;
assign img[ 4293] = 221;
assign img[ 4294] = 253;
assign img[ 4295] = 255;
assign img[ 4296] = 255;
assign img[ 4297] = 255;
assign img[ 4298] = 255;
assign img[ 4299] = 255;
assign img[ 4300] = 255;
assign img[ 4301] = 255;
assign img[ 4302] = 255;
assign img[ 4303] = 255;
assign img[ 4304] = 255;
assign img[ 4305] = 255;
assign img[ 4306] = 255;
assign img[ 4307] = 255;
assign img[ 4308] = 255;
assign img[ 4309] = 255;
assign img[ 4310] = 238;
assign img[ 4311] = 238;
assign img[ 4312] = 254;
assign img[ 4313] = 255;
assign img[ 4314] = 255;
assign img[ 4315] = 255;
assign img[ 4316] = 255;
assign img[ 4317] = 255;
assign img[ 4318] = 255;
assign img[ 4319] = 159;
assign img[ 4320] = 137;
assign img[ 4321] = 238;
assign img[ 4322] = 254;
assign img[ 4323] = 255;
assign img[ 4324] = 255;
assign img[ 4325] = 223;
assign img[ 4326] = 221;
assign img[ 4327] = 221;
assign img[ 4328] = 253;
assign img[ 4329] = 223;
assign img[ 4330] = 253;
assign img[ 4331] = 255;
assign img[ 4332] = 239;
assign img[ 4333] = 238;
assign img[ 4334] = 238;
assign img[ 4335] = 174;
assign img[ 4336] = 250;
assign img[ 4337] = 171;
assign img[ 4338] = 234;
assign img[ 4339] = 254;
assign img[ 4340] = 221;
assign img[ 4341] = 221;
assign img[ 4342] = 253;
assign img[ 4343] = 255;
assign img[ 4344] = 255;
assign img[ 4345] = 255;
assign img[ 4346] = 238;
assign img[ 4347] = 238;
assign img[ 4348] = 238;
assign img[ 4349] = 238;
assign img[ 4350] = 238;
assign img[ 4351] = 255;
assign img[ 4352] = 96;
assign img[ 4353] = 238;
assign img[ 4354] = 254;
assign img[ 4355] = 207;
assign img[ 4356] = 140;
assign img[ 4357] = 136;
assign img[ 4358] = 136;
assign img[ 4359] = 236;
assign img[ 4360] = 238;
assign img[ 4361] = 255;
assign img[ 4362] = 238;
assign img[ 4363] = 254;
assign img[ 4364] = 239;
assign img[ 4365] = 255;
assign img[ 4366] = 239;
assign img[ 4367] = 238;
assign img[ 4368] = 238;
assign img[ 4369] = 238;
assign img[ 4370] = 238;
assign img[ 4371] = 238;
assign img[ 4372] = 238;
assign img[ 4373] = 238;
assign img[ 4374] = 238;
assign img[ 4375] = 238;
assign img[ 4376] = 238;
assign img[ 4377] = 238;
assign img[ 4378] = 238;
assign img[ 4379] = 238;
assign img[ 4380] = 206;
assign img[ 4381] = 255;
assign img[ 4382] = 223;
assign img[ 4383] = 221;
assign img[ 4384] = 221;
assign img[ 4385] = 253;
assign img[ 4386] = 255;
assign img[ 4387] = 255;
assign img[ 4388] = 255;
assign img[ 4389] = 239;
assign img[ 4390] = 254;
assign img[ 4391] = 255;
assign img[ 4392] = 255;
assign img[ 4393] = 255;
assign img[ 4394] = 255;
assign img[ 4395] = 255;
assign img[ 4396] = 238;
assign img[ 4397] = 238;
assign img[ 4398] = 238;
assign img[ 4399] = 206;
assign img[ 4400] = 254;
assign img[ 4401] = 255;
assign img[ 4402] = 239;
assign img[ 4403] = 238;
assign img[ 4404] = 238;
assign img[ 4405] = 238;
assign img[ 4406] = 238;
assign img[ 4407] = 238;
assign img[ 4408] = 238;
assign img[ 4409] = 238;
assign img[ 4410] = 206;
assign img[ 4411] = 204;
assign img[ 4412] = 236;
assign img[ 4413] = 174;
assign img[ 4414] = 238;
assign img[ 4415] = 254;
assign img[ 4416] = 238;
assign img[ 4417] = 255;
assign img[ 4418] = 255;
assign img[ 4419] = 255;
assign img[ 4420] = 255;
assign img[ 4421] = 223;
assign img[ 4422] = 253;
assign img[ 4423] = 255;
assign img[ 4424] = 238;
assign img[ 4425] = 238;
assign img[ 4426] = 254;
assign img[ 4427] = 255;
assign img[ 4428] = 255;
assign img[ 4429] = 255;
assign img[ 4430] = 238;
assign img[ 4431] = 255;
assign img[ 4432] = 223;
assign img[ 4433] = 255;
assign img[ 4434] = 255;
assign img[ 4435] = 255;
assign img[ 4436] = 255;
assign img[ 4437] = 255;
assign img[ 4438] = 255;
assign img[ 4439] = 255;
assign img[ 4440] = 191;
assign img[ 4441] = 255;
assign img[ 4442] = 255;
assign img[ 4443] = 255;
assign img[ 4444] = 255;
assign img[ 4445] = 255;
assign img[ 4446] = 255;
assign img[ 4447] = 239;
assign img[ 4448] = 204;
assign img[ 4449] = 204;
assign img[ 4450] = 252;
assign img[ 4451] = 223;
assign img[ 4452] = 253;
assign img[ 4453] = 239;
assign img[ 4454] = 204;
assign img[ 4455] = 236;
assign img[ 4456] = 238;
assign img[ 4457] = 255;
assign img[ 4458] = 255;
assign img[ 4459] = 255;
assign img[ 4460] = 255;
assign img[ 4461] = 255;
assign img[ 4462] = 255;
assign img[ 4463] = 255;
assign img[ 4464] = 255;
assign img[ 4465] = 255;
assign img[ 4466] = 255;
assign img[ 4467] = 255;
assign img[ 4468] = 255;
assign img[ 4469] = 239;
assign img[ 4470] = 238;
assign img[ 4471] = 238;
assign img[ 4472] = 238;
assign img[ 4473] = 239;
assign img[ 4474] = 238;
assign img[ 4475] = 174;
assign img[ 4476] = 200;
assign img[ 4477] = 252;
assign img[ 4478] = 255;
assign img[ 4479] = 255;
assign img[ 4480] = 96;
assign img[ 4481] = 223;
assign img[ 4482] = 253;
assign img[ 4483] = 207;
assign img[ 4484] = 204;
assign img[ 4485] = 204;
assign img[ 4486] = 204;
assign img[ 4487] = 236;
assign img[ 4488] = 238;
assign img[ 4489] = 238;
assign img[ 4490] = 238;
assign img[ 4491] = 238;
assign img[ 4492] = 238;
assign img[ 4493] = 238;
assign img[ 4494] = 238;
assign img[ 4495] = 206;
assign img[ 4496] = 220;
assign img[ 4497] = 221;
assign img[ 4498] = 221;
assign img[ 4499] = 205;
assign img[ 4500] = 220;
assign img[ 4501] = 253;
assign img[ 4502] = 255;
assign img[ 4503] = 255;
assign img[ 4504] = 255;
assign img[ 4505] = 255;
assign img[ 4506] = 223;
assign img[ 4507] = 255;
assign img[ 4508] = 223;
assign img[ 4509] = 255;
assign img[ 4510] = 239;
assign img[ 4511] = 190;
assign img[ 4512] = 139;
assign img[ 4513] = 238;
assign img[ 4514] = 238;
assign img[ 4515] = 238;
assign img[ 4516] = 238;
assign img[ 4517] = 238;
assign img[ 4518] = 238;
assign img[ 4519] = 238;
assign img[ 4520] = 238;
assign img[ 4521] = 238;
assign img[ 4522] = 238;
assign img[ 4523] = 254;
assign img[ 4524] = 254;
assign img[ 4525] = 255;
assign img[ 4526] = 255;
assign img[ 4527] = 255;
assign img[ 4528] = 255;
assign img[ 4529] = 255;
assign img[ 4530] = 255;
assign img[ 4531] = 255;
assign img[ 4532] = 255;
assign img[ 4533] = 255;
assign img[ 4534] = 255;
assign img[ 4535] = 255;
assign img[ 4536] = 255;
assign img[ 4537] = 255;
assign img[ 4538] = 255;
assign img[ 4539] = 255;
assign img[ 4540] = 255;
assign img[ 4541] = 223;
assign img[ 4542] = 255;
assign img[ 4543] = 255;
assign img[ 4544] = 255;
assign img[ 4545] = 255;
assign img[ 4546] = 223;
assign img[ 4547] = 255;
assign img[ 4548] = 255;
assign img[ 4549] = 255;
assign img[ 4550] = 255;
assign img[ 4551] = 255;
assign img[ 4552] = 255;
assign img[ 4553] = 255;
assign img[ 4554] = 255;
assign img[ 4555] = 255;
assign img[ 4556] = 255;
assign img[ 4557] = 239;
assign img[ 4558] = 238;
assign img[ 4559] = 255;
assign img[ 4560] = 223;
assign img[ 4561] = 255;
assign img[ 4562] = 255;
assign img[ 4563] = 255;
assign img[ 4564] = 255;
assign img[ 4565] = 255;
assign img[ 4566] = 255;
assign img[ 4567] = 255;
assign img[ 4568] = 223;
assign img[ 4569] = 255;
assign img[ 4570] = 239;
assign img[ 4571] = 239;
assign img[ 4572] = 238;
assign img[ 4573] = 238;
assign img[ 4574] = 238;
assign img[ 4575] = 223;
assign img[ 4576] = 236;
assign img[ 4577] = 239;
assign img[ 4578] = 238;
assign img[ 4579] = 238;
assign img[ 4580] = 238;
assign img[ 4581] = 255;
assign img[ 4582] = 255;
assign img[ 4583] = 255;
assign img[ 4584] = 255;
assign img[ 4585] = 255;
assign img[ 4586] = 255;
assign img[ 4587] = 255;
assign img[ 4588] = 221;
assign img[ 4589] = 205;
assign img[ 4590] = 236;
assign img[ 4591] = 238;
assign img[ 4592] = 138;
assign img[ 4593] = 236;
assign img[ 4594] = 238;
assign img[ 4595] = 255;
assign img[ 4596] = 255;
assign img[ 4597] = 255;
assign img[ 4598] = 238;
assign img[ 4599] = 238;
assign img[ 4600] = 238;
assign img[ 4601] = 255;
assign img[ 4602] = 239;
assign img[ 4603] = 238;
assign img[ 4604] = 238;
assign img[ 4605] = 255;
assign img[ 4606] = 254;
assign img[ 4607] = 255;
assign img[ 4608] = 96;
assign img[ 4609] = 207;
assign img[ 4610] = 253;
assign img[ 4611] = 255;
assign img[ 4612] = 223;
assign img[ 4613] = 221;
assign img[ 4614] = 253;
assign img[ 4615] = 239;
assign img[ 4616] = 238;
assign img[ 4617] = 238;
assign img[ 4618] = 238;
assign img[ 4619] = 238;
assign img[ 4620] = 204;
assign img[ 4621] = 204;
assign img[ 4622] = 253;
assign img[ 4623] = 207;
assign img[ 4624] = 204;
assign img[ 4625] = 236;
assign img[ 4626] = 238;
assign img[ 4627] = 206;
assign img[ 4628] = 220;
assign img[ 4629] = 253;
assign img[ 4630] = 255;
assign img[ 4631] = 255;
assign img[ 4632] = 255;
assign img[ 4633] = 255;
assign img[ 4634] = 204;
assign img[ 4635] = 238;
assign img[ 4636] = 238;
assign img[ 4637] = 255;
assign img[ 4638] = 239;
assign img[ 4639] = 174;
assign img[ 4640] = 170;
assign img[ 4641] = 238;
assign img[ 4642] = 238;
assign img[ 4643] = 238;
assign img[ 4644] = 238;
assign img[ 4645] = 255;
assign img[ 4646] = 255;
assign img[ 4647] = 255;
assign img[ 4648] = 238;
assign img[ 4649] = 238;
assign img[ 4650] = 222;
assign img[ 4651] = 255;
assign img[ 4652] = 255;
assign img[ 4653] = 255;
assign img[ 4654] = 255;
assign img[ 4655] = 255;
assign img[ 4656] = 255;
assign img[ 4657] = 255;
assign img[ 4658] = 255;
assign img[ 4659] = 255;
assign img[ 4660] = 255;
assign img[ 4661] = 255;
assign img[ 4662] = 255;
assign img[ 4663] = 255;
assign img[ 4664] = 255;
assign img[ 4665] = 255;
assign img[ 4666] = 223;
assign img[ 4667] = 255;
assign img[ 4668] = 223;
assign img[ 4669] = 157;
assign img[ 4670] = 249;
assign img[ 4671] = 255;
assign img[ 4672] = 255;
assign img[ 4673] = 255;
assign img[ 4674] = 191;
assign img[ 4675] = 139;
assign img[ 4676] = 232;
assign img[ 4677] = 206;
assign img[ 4678] = 236;
assign img[ 4679] = 238;
assign img[ 4680] = 238;
assign img[ 4681] = 254;
assign img[ 4682] = 254;
assign img[ 4683] = 238;
assign img[ 4684] = 238;
assign img[ 4685] = 238;
assign img[ 4686] = 238;
assign img[ 4687] = 255;
assign img[ 4688] = 255;
assign img[ 4689] = 255;
assign img[ 4690] = 223;
assign img[ 4691] = 255;
assign img[ 4692] = 255;
assign img[ 4693] = 255;
assign img[ 4694] = 255;
assign img[ 4695] = 255;
assign img[ 4696] = 223;
assign img[ 4697] = 255;
assign img[ 4698] = 255;
assign img[ 4699] = 255;
assign img[ 4700] = 255;
assign img[ 4701] = 239;
assign img[ 4702] = 238;
assign img[ 4703] = 206;
assign img[ 4704] = 156;
assign img[ 4705] = 153;
assign img[ 4706] = 249;
assign img[ 4707] = 255;
assign img[ 4708] = 255;
assign img[ 4709] = 255;
assign img[ 4710] = 206;
assign img[ 4711] = 204;
assign img[ 4712] = 238;
assign img[ 4713] = 238;
assign img[ 4714] = 238;
assign img[ 4715] = 238;
assign img[ 4716] = 238;
assign img[ 4717] = 255;
assign img[ 4718] = 255;
assign img[ 4719] = 255;
assign img[ 4720] = 255;
assign img[ 4721] = 255;
assign img[ 4722] = 255;
assign img[ 4723] = 255;
assign img[ 4724] = 221;
assign img[ 4725] = 253;
assign img[ 4726] = 238;
assign img[ 4727] = 238;
assign img[ 4728] = 255;
assign img[ 4729] = 255;
assign img[ 4730] = 187;
assign img[ 4731] = 223;
assign img[ 4732] = 221;
assign img[ 4733] = 255;
assign img[ 4734] = 223;
assign img[ 4735] = 253;
assign img[ 4736] = 96;
assign img[ 4737] = 238;
assign img[ 4738] = 238;
assign img[ 4739] = 223;
assign img[ 4740] = 253;
assign img[ 4741] = 238;
assign img[ 4742] = 255;
assign img[ 4743] = 255;
assign img[ 4744] = 255;
assign img[ 4745] = 255;
assign img[ 4746] = 255;
assign img[ 4747] = 239;
assign img[ 4748] = 254;
assign img[ 4749] = 255;
assign img[ 4750] = 255;
assign img[ 4751] = 223;
assign img[ 4752] = 205;
assign img[ 4753] = 238;
assign img[ 4754] = 238;
assign img[ 4755] = 174;
assign img[ 4756] = 170;
assign img[ 4757] = 238;
assign img[ 4758] = 238;
assign img[ 4759] = 238;
assign img[ 4760] = 254;
assign img[ 4761] = 255;
assign img[ 4762] = 239;
assign img[ 4763] = 238;
assign img[ 4764] = 238;
assign img[ 4765] = 238;
assign img[ 4766] = 238;
assign img[ 4767] = 238;
assign img[ 4768] = 254;
assign img[ 4769] = 255;
assign img[ 4770] = 255;
assign img[ 4771] = 255;
assign img[ 4772] = 255;
assign img[ 4773] = 255;
assign img[ 4774] = 255;
assign img[ 4775] = 239;
assign img[ 4776] = 238;
assign img[ 4777] = 238;
assign img[ 4778] = 254;
assign img[ 4779] = 223;
assign img[ 4780] = 253;
assign img[ 4781] = 255;
assign img[ 4782] = 255;
assign img[ 4783] = 255;
assign img[ 4784] = 255;
assign img[ 4785] = 255;
assign img[ 4786] = 255;
assign img[ 4787] = 255;
assign img[ 4788] = 255;
assign img[ 4789] = 255;
assign img[ 4790] = 255;
assign img[ 4791] = 255;
assign img[ 4792] = 255;
assign img[ 4793] = 255;
assign img[ 4794] = 254;
assign img[ 4795] = 255;
assign img[ 4796] = 255;
assign img[ 4797] = 223;
assign img[ 4798] = 255;
assign img[ 4799] = 255;
assign img[ 4800] = 255;
assign img[ 4801] = 255;
assign img[ 4802] = 223;
assign img[ 4803] = 255;
assign img[ 4804] = 255;
assign img[ 4805] = 223;
assign img[ 4806] = 253;
assign img[ 4807] = 239;
assign img[ 4808] = 238;
assign img[ 4809] = 238;
assign img[ 4810] = 238;
assign img[ 4811] = 255;
assign img[ 4812] = 255;
assign img[ 4813] = 238;
assign img[ 4814] = 254;
assign img[ 4815] = 255;
assign img[ 4816] = 255;
assign img[ 4817] = 255;
assign img[ 4818] = 255;
assign img[ 4819] = 255;
assign img[ 4820] = 223;
assign img[ 4821] = 221;
assign img[ 4822] = 255;
assign img[ 4823] = 255;
assign img[ 4824] = 255;
assign img[ 4825] = 255;
assign img[ 4826] = 255;
assign img[ 4827] = 255;
assign img[ 4828] = 255;
assign img[ 4829] = 255;
assign img[ 4830] = 255;
assign img[ 4831] = 255;
assign img[ 4832] = 255;
assign img[ 4833] = 238;
assign img[ 4834] = 238;
assign img[ 4835] = 255;
assign img[ 4836] = 255;
assign img[ 4837] = 239;
assign img[ 4838] = 174;
assign img[ 4839] = 170;
assign img[ 4840] = 234;
assign img[ 4841] = 239;
assign img[ 4842] = 238;
assign img[ 4843] = 239;
assign img[ 4844] = 255;
assign img[ 4845] = 255;
assign img[ 4846] = 255;
assign img[ 4847] = 255;
assign img[ 4848] = 238;
assign img[ 4849] = 238;
assign img[ 4850] = 238;
assign img[ 4851] = 238;
assign img[ 4852] = 238;
assign img[ 4853] = 238;
assign img[ 4854] = 238;
assign img[ 4855] = 255;
assign img[ 4856] = 238;
assign img[ 4857] = 255;
assign img[ 4858] = 255;
assign img[ 4859] = 255;
assign img[ 4860] = 238;
assign img[ 4861] = 238;
assign img[ 4862] = 238;
assign img[ 4863] = 238;
assign img[ 4864] = 96;
assign img[ 4865] = 239;
assign img[ 4866] = 238;
assign img[ 4867] = 238;
assign img[ 4868] = 238;
assign img[ 4869] = 238;
assign img[ 4870] = 206;
assign img[ 4871] = 254;
assign img[ 4872] = 255;
assign img[ 4873] = 254;
assign img[ 4874] = 255;
assign img[ 4875] = 238;
assign img[ 4876] = 238;
assign img[ 4877] = 254;
assign img[ 4878] = 255;
assign img[ 4879] = 239;
assign img[ 4880] = 238;
assign img[ 4881] = 239;
assign img[ 4882] = 238;
assign img[ 4883] = 222;
assign img[ 4884] = 204;
assign img[ 4885] = 253;
assign img[ 4886] = 255;
assign img[ 4887] = 255;
assign img[ 4888] = 255;
assign img[ 4889] = 239;
assign img[ 4890] = 204;
assign img[ 4891] = 236;
assign img[ 4892] = 238;
assign img[ 4893] = 255;
assign img[ 4894] = 255;
assign img[ 4895] = 207;
assign img[ 4896] = 204;
assign img[ 4897] = 236;
assign img[ 4898] = 238;
assign img[ 4899] = 238;
assign img[ 4900] = 238;
assign img[ 4901] = 238;
assign img[ 4902] = 254;
assign img[ 4903] = 255;
assign img[ 4904] = 255;
assign img[ 4905] = 255;
assign img[ 4906] = 255;
assign img[ 4907] = 223;
assign img[ 4908] = 221;
assign img[ 4909] = 221;
assign img[ 4910] = 253;
assign img[ 4911] = 255;
assign img[ 4912] = 255;
assign img[ 4913] = 255;
assign img[ 4914] = 255;
assign img[ 4915] = 255;
assign img[ 4916] = 255;
assign img[ 4917] = 255;
assign img[ 4918] = 255;
assign img[ 4919] = 255;
assign img[ 4920] = 255;
assign img[ 4921] = 255;
assign img[ 4922] = 239;
assign img[ 4923] = 238;
assign img[ 4924] = 238;
assign img[ 4925] = 255;
assign img[ 4926] = 238;
assign img[ 4927] = 255;
assign img[ 4928] = 255;
assign img[ 4929] = 255;
assign img[ 4930] = 255;
assign img[ 4931] = 255;
assign img[ 4932] = 255;
assign img[ 4933] = 255;
assign img[ 4934] = 238;
assign img[ 4935] = 238;
assign img[ 4936] = 238;
assign img[ 4937] = 255;
assign img[ 4938] = 255;
assign img[ 4939] = 255;
assign img[ 4940] = 255;
assign img[ 4941] = 255;
assign img[ 4942] = 255;
assign img[ 4943] = 255;
assign img[ 4944] = 255;
assign img[ 4945] = 255;
assign img[ 4946] = 223;
assign img[ 4947] = 221;
assign img[ 4948] = 221;
assign img[ 4949] = 221;
assign img[ 4950] = 253;
assign img[ 4951] = 255;
assign img[ 4952] = 255;
assign img[ 4953] = 255;
assign img[ 4954] = 239;
assign img[ 4955] = 239;
assign img[ 4956] = 238;
assign img[ 4957] = 238;
assign img[ 4958] = 238;
assign img[ 4959] = 223;
assign img[ 4960] = 253;
assign img[ 4961] = 239;
assign img[ 4962] = 254;
assign img[ 4963] = 255;
assign img[ 4964] = 255;
assign img[ 4965] = 223;
assign img[ 4966] = 221;
assign img[ 4967] = 221;
assign img[ 4968] = 253;
assign img[ 4969] = 255;
assign img[ 4970] = 255;
assign img[ 4971] = 223;
assign img[ 4972] = 221;
assign img[ 4973] = 221;
assign img[ 4974] = 236;
assign img[ 4975] = 238;
assign img[ 4976] = 238;
assign img[ 4977] = 238;
assign img[ 4978] = 206;
assign img[ 4979] = 204;
assign img[ 4980] = 236;
assign img[ 4981] = 238;
assign img[ 4982] = 238;
assign img[ 4983] = 238;
assign img[ 4984] = 238;
assign img[ 4985] = 255;
assign img[ 4986] = 238;
assign img[ 4987] = 239;
assign img[ 4988] = 255;
assign img[ 4989] = 255;
assign img[ 4990] = 239;
assign img[ 4991] = 238;
assign img[ 4992] = 96;
assign img[ 4993] = 255;
assign img[ 4994] = 255;
assign img[ 4995] = 207;
assign img[ 4996] = 204;
assign img[ 4997] = 204;
assign img[ 4998] = 204;
assign img[ 4999] = 236;
assign img[ 5000] = 238;
assign img[ 5001] = 255;
assign img[ 5002] = 255;
assign img[ 5003] = 255;
assign img[ 5004] = 255;
assign img[ 5005] = 255;
assign img[ 5006] = 223;
assign img[ 5007] = 255;
assign img[ 5008] = 223;
assign img[ 5009] = 221;
assign img[ 5010] = 236;
assign img[ 5011] = 255;
assign img[ 5012] = 255;
assign img[ 5013] = 255;
assign img[ 5014] = 239;
assign img[ 5015] = 255;
assign img[ 5016] = 255;
assign img[ 5017] = 255;
assign img[ 5018] = 221;
assign img[ 5019] = 253;
assign img[ 5020] = 255;
assign img[ 5021] = 255;
assign img[ 5022] = 255;
assign img[ 5023] = 223;
assign img[ 5024] = 221;
assign img[ 5025] = 255;
assign img[ 5026] = 255;
assign img[ 5027] = 255;
assign img[ 5028] = 255;
assign img[ 5029] = 255;
assign img[ 5030] = 255;
assign img[ 5031] = 255;
assign img[ 5032] = 255;
assign img[ 5033] = 255;
assign img[ 5034] = 255;
assign img[ 5035] = 255;
assign img[ 5036] = 255;
assign img[ 5037] = 255;
assign img[ 5038] = 255;
assign img[ 5039] = 255;
assign img[ 5040] = 255;
assign img[ 5041] = 255;
assign img[ 5042] = 255;
assign img[ 5043] = 255;
assign img[ 5044] = 255;
assign img[ 5045] = 255;
assign img[ 5046] = 255;
assign img[ 5047] = 255;
assign img[ 5048] = 255;
assign img[ 5049] = 255;
assign img[ 5050] = 239;
assign img[ 5051] = 238;
assign img[ 5052] = 238;
assign img[ 5053] = 207;
assign img[ 5054] = 238;
assign img[ 5055] = 254;
assign img[ 5056] = 255;
assign img[ 5057] = 255;
assign img[ 5058] = 238;
assign img[ 5059] = 238;
assign img[ 5060] = 238;
assign img[ 5061] = 239;
assign img[ 5062] = 238;
assign img[ 5063] = 238;
assign img[ 5064] = 238;
assign img[ 5065] = 238;
assign img[ 5066] = 254;
assign img[ 5067] = 255;
assign img[ 5068] = 255;
assign img[ 5069] = 239;
assign img[ 5070] = 238;
assign img[ 5071] = 255;
assign img[ 5072] = 239;
assign img[ 5073] = 238;
assign img[ 5074] = 238;
assign img[ 5075] = 238;
assign img[ 5076] = 238;
assign img[ 5077] = 238;
assign img[ 5078] = 238;
assign img[ 5079] = 238;
assign img[ 5080] = 238;
assign img[ 5081] = 255;
assign img[ 5082] = 255;
assign img[ 5083] = 223;
assign img[ 5084] = 253;
assign img[ 5085] = 255;
assign img[ 5086] = 255;
assign img[ 5087] = 191;
assign img[ 5088] = 139;
assign img[ 5089] = 206;
assign img[ 5090] = 238;
assign img[ 5091] = 238;
assign img[ 5092] = 238;
assign img[ 5093] = 238;
assign img[ 5094] = 204;
assign img[ 5095] = 236;
assign img[ 5096] = 254;
assign img[ 5097] = 255;
assign img[ 5098] = 238;
assign img[ 5099] = 238;
assign img[ 5100] = 254;
assign img[ 5101] = 255;
assign img[ 5102] = 255;
assign img[ 5103] = 255;
assign img[ 5104] = 255;
assign img[ 5105] = 239;
assign img[ 5106] = 238;
assign img[ 5107] = 238;
assign img[ 5108] = 238;
assign img[ 5109] = 238;
assign img[ 5110] = 254;
assign img[ 5111] = 255;
assign img[ 5112] = 255;
assign img[ 5113] = 255;
assign img[ 5114] = 204;
assign img[ 5115] = 236;
assign img[ 5116] = 206;
assign img[ 5117] = 252;
assign img[ 5118] = 255;
assign img[ 5119] = 255;
assign img[ 5120] = 96;
assign img[ 5121] = 238;
assign img[ 5122] = 238;
assign img[ 5123] = 238;
assign img[ 5124] = 254;
assign img[ 5125] = 255;
assign img[ 5126] = 255;
assign img[ 5127] = 255;
assign img[ 5128] = 255;
assign img[ 5129] = 255;
assign img[ 5130] = 255;
assign img[ 5131] = 223;
assign img[ 5132] = 204;
assign img[ 5133] = 221;
assign img[ 5134] = 221;
assign img[ 5135] = 157;
assign img[ 5136] = 221;
assign img[ 5137] = 253;
assign img[ 5138] = 255;
assign img[ 5139] = 207;
assign img[ 5140] = 254;
assign img[ 5141] = 255;
assign img[ 5142] = 223;
assign img[ 5143] = 255;
assign img[ 5144] = 255;
assign img[ 5145] = 255;
assign img[ 5146] = 239;
assign img[ 5147] = 238;
assign img[ 5148] = 238;
assign img[ 5149] = 238;
assign img[ 5150] = 238;
assign img[ 5151] = 174;
assign img[ 5152] = 187;
assign img[ 5153] = 251;
assign img[ 5154] = 255;
assign img[ 5155] = 255;
assign img[ 5156] = 255;
assign img[ 5157] = 255;
assign img[ 5158] = 255;
assign img[ 5159] = 255;
assign img[ 5160] = 255;
assign img[ 5161] = 255;
assign img[ 5162] = 255;
assign img[ 5163] = 255;
assign img[ 5164] = 255;
assign img[ 5165] = 239;
assign img[ 5166] = 238;
assign img[ 5167] = 255;
assign img[ 5168] = 255;
assign img[ 5169] = 255;
assign img[ 5170] = 255;
assign img[ 5171] = 255;
assign img[ 5172] = 255;
assign img[ 5173] = 255;
assign img[ 5174] = 255;
assign img[ 5175] = 255;
assign img[ 5176] = 255;
assign img[ 5177] = 255;
assign img[ 5178] = 239;
assign img[ 5179] = 255;
assign img[ 5180] = 255;
assign img[ 5181] = 207;
assign img[ 5182] = 204;
assign img[ 5183] = 238;
assign img[ 5184] = 238;
assign img[ 5185] = 238;
assign img[ 5186] = 238;
assign img[ 5187] = 238;
assign img[ 5188] = 206;
assign img[ 5189] = 205;
assign img[ 5190] = 253;
assign img[ 5191] = 255;
assign img[ 5192] = 255;
assign img[ 5193] = 255;
assign img[ 5194] = 255;
assign img[ 5195] = 255;
assign img[ 5196] = 238;
assign img[ 5197] = 255;
assign img[ 5198] = 254;
assign img[ 5199] = 255;
assign img[ 5200] = 207;
assign img[ 5201] = 238;
assign img[ 5202] = 238;
assign img[ 5203] = 238;
assign img[ 5204] = 238;
assign img[ 5205] = 238;
assign img[ 5206] = 238;
assign img[ 5207] = 238;
assign img[ 5208] = 238;
assign img[ 5209] = 255;
assign img[ 5210] = 255;
assign img[ 5211] = 255;
assign img[ 5212] = 255;
assign img[ 5213] = 255;
assign img[ 5214] = 255;
assign img[ 5215] = 191;
assign img[ 5216] = 255;
assign img[ 5217] = 255;
assign img[ 5218] = 238;
assign img[ 5219] = 238;
assign img[ 5220] = 254;
assign img[ 5221] = 255;
assign img[ 5222] = 191;
assign img[ 5223] = 187;
assign img[ 5224] = 251;
assign img[ 5225] = 255;
assign img[ 5226] = 255;
assign img[ 5227] = 255;
assign img[ 5228] = 255;
assign img[ 5229] = 255;
assign img[ 5230] = 255;
assign img[ 5231] = 255;
assign img[ 5232] = 140;
assign img[ 5233] = 152;
assign img[ 5234] = 152;
assign img[ 5235] = 221;
assign img[ 5236] = 205;
assign img[ 5237] = 236;
assign img[ 5238] = 238;
assign img[ 5239] = 238;
assign img[ 5240] = 238;
assign img[ 5241] = 238;
assign img[ 5242] = 170;
assign img[ 5243] = 238;
assign img[ 5244] = 220;
assign img[ 5245] = 255;
assign img[ 5246] = 255;
assign img[ 5247] = 255;
assign img[ 5248] = 96;
assign img[ 5249] = 206;
assign img[ 5250] = 220;
assign img[ 5251] = 253;
assign img[ 5252] = 255;
assign img[ 5253] = 223;
assign img[ 5254] = 221;
assign img[ 5255] = 253;
assign img[ 5256] = 255;
assign img[ 5257] = 255;
assign img[ 5258] = 255;
assign img[ 5259] = 223;
assign img[ 5260] = 221;
assign img[ 5261] = 221;
assign img[ 5262] = 205;
assign img[ 5263] = 206;
assign img[ 5264] = 238;
assign img[ 5265] = 255;
assign img[ 5266] = 255;
assign img[ 5267] = 239;
assign img[ 5268] = 238;
assign img[ 5269] = 238;
assign img[ 5270] = 238;
assign img[ 5271] = 238;
assign img[ 5272] = 254;
assign img[ 5273] = 255;
assign img[ 5274] = 255;
assign img[ 5275] = 255;
assign img[ 5276] = 255;
assign img[ 5277] = 255;
assign img[ 5278] = 239;
assign img[ 5279] = 223;
assign img[ 5280] = 157;
assign img[ 5281] = 255;
assign img[ 5282] = 255;
assign img[ 5283] = 255;
assign img[ 5284] = 255;
assign img[ 5285] = 255;
assign img[ 5286] = 255;
assign img[ 5287] = 239;
assign img[ 5288] = 238;
assign img[ 5289] = 206;
assign img[ 5290] = 238;
assign img[ 5291] = 238;
assign img[ 5292] = 238;
assign img[ 5293] = 255;
assign img[ 5294] = 255;
assign img[ 5295] = 255;
assign img[ 5296] = 255;
assign img[ 5297] = 255;
assign img[ 5298] = 255;
assign img[ 5299] = 223;
assign img[ 5300] = 221;
assign img[ 5301] = 255;
assign img[ 5302] = 255;
assign img[ 5303] = 255;
assign img[ 5304] = 255;
assign img[ 5305] = 255;
assign img[ 5306] = 239;
assign img[ 5307] = 238;
assign img[ 5308] = 238;
assign img[ 5309] = 238;
assign img[ 5310] = 238;
assign img[ 5311] = 254;
assign img[ 5312] = 255;
assign img[ 5313] = 255;
assign img[ 5314] = 255;
assign img[ 5315] = 255;
assign img[ 5316] = 255;
assign img[ 5317] = 255;
assign img[ 5318] = 238;
assign img[ 5319] = 238;
assign img[ 5320] = 238;
assign img[ 5321] = 254;
assign img[ 5322] = 255;
assign img[ 5323] = 255;
assign img[ 5324] = 255;
assign img[ 5325] = 255;
assign img[ 5326] = 255;
assign img[ 5327] = 255;
assign img[ 5328] = 255;
assign img[ 5329] = 255;
assign img[ 5330] = 255;
assign img[ 5331] = 255;
assign img[ 5332] = 238;
assign img[ 5333] = 255;
assign img[ 5334] = 223;
assign img[ 5335] = 255;
assign img[ 5336] = 255;
assign img[ 5337] = 255;
assign img[ 5338] = 239;
assign img[ 5339] = 238;
assign img[ 5340] = 238;
assign img[ 5341] = 238;
assign img[ 5342] = 254;
assign img[ 5343] = 191;
assign img[ 5344] = 223;
assign img[ 5345] = 205;
assign img[ 5346] = 252;
assign img[ 5347] = 255;
assign img[ 5348] = 255;
assign img[ 5349] = 255;
assign img[ 5350] = 239;
assign img[ 5351] = 238;
assign img[ 5352] = 238;
assign img[ 5353] = 255;
assign img[ 5354] = 255;
assign img[ 5355] = 255;
assign img[ 5356] = 255;
assign img[ 5357] = 255;
assign img[ 5358] = 255;
assign img[ 5359] = 255;
assign img[ 5360] = 255;
assign img[ 5361] = 255;
assign img[ 5362] = 255;
assign img[ 5363] = 223;
assign img[ 5364] = 221;
assign img[ 5365] = 253;
assign img[ 5366] = 255;
assign img[ 5367] = 255;
assign img[ 5368] = 255;
assign img[ 5369] = 223;
assign img[ 5370] = 221;
assign img[ 5371] = 205;
assign img[ 5372] = 236;
assign img[ 5373] = 238;
assign img[ 5374] = 204;
assign img[ 5375] = 236;
assign img[ 5376] = 96;
assign img[ 5377] = 238;
assign img[ 5378] = 254;
assign img[ 5379] = 223;
assign img[ 5380] = 221;
assign img[ 5381] = 221;
assign img[ 5382] = 253;
assign img[ 5383] = 239;
assign img[ 5384] = 238;
assign img[ 5385] = 239;
assign img[ 5386] = 206;
assign img[ 5387] = 204;
assign img[ 5388] = 236;
assign img[ 5389] = 238;
assign img[ 5390] = 238;
assign img[ 5391] = 238;
assign img[ 5392] = 238;
assign img[ 5393] = 238;
assign img[ 5394] = 238;
assign img[ 5395] = 238;
assign img[ 5396] = 238;
assign img[ 5397] = 238;
assign img[ 5398] = 238;
assign img[ 5399] = 238;
assign img[ 5400] = 238;
assign img[ 5401] = 255;
assign img[ 5402] = 207;
assign img[ 5403] = 238;
assign img[ 5404] = 238;
assign img[ 5405] = 255;
assign img[ 5406] = 223;
assign img[ 5407] = 221;
assign img[ 5408] = 221;
assign img[ 5409] = 253;
assign img[ 5410] = 255;
assign img[ 5411] = 255;
assign img[ 5412] = 223;
assign img[ 5413] = 221;
assign img[ 5414] = 253;
assign img[ 5415] = 255;
assign img[ 5416] = 238;
assign img[ 5417] = 238;
assign img[ 5418] = 255;
assign img[ 5419] = 255;
assign img[ 5420] = 254;
assign img[ 5421] = 255;
assign img[ 5422] = 238;
assign img[ 5423] = 239;
assign img[ 5424] = 238;
assign img[ 5425] = 238;
assign img[ 5426] = 238;
assign img[ 5427] = 223;
assign img[ 5428] = 206;
assign img[ 5429] = 255;
assign img[ 5430] = 255;
assign img[ 5431] = 255;
assign img[ 5432] = 239;
assign img[ 5433] = 238;
assign img[ 5434] = 238;
assign img[ 5435] = 238;
assign img[ 5436] = 238;
assign img[ 5437] = 255;
assign img[ 5438] = 255;
assign img[ 5439] = 255;
assign img[ 5440] = 255;
assign img[ 5441] = 255;
assign img[ 5442] = 223;
assign img[ 5443] = 255;
assign img[ 5444] = 255;
assign img[ 5445] = 255;
assign img[ 5446] = 255;
assign img[ 5447] = 255;
assign img[ 5448] = 238;
assign img[ 5449] = 238;
assign img[ 5450] = 254;
assign img[ 5451] = 255;
assign img[ 5452] = 239;
assign img[ 5453] = 238;
assign img[ 5454] = 238;
assign img[ 5455] = 238;
assign img[ 5456] = 238;
assign img[ 5457] = 238;
assign img[ 5458] = 238;
assign img[ 5459] = 238;
assign img[ 5460] = 254;
assign img[ 5461] = 239;
assign img[ 5462] = 238;
assign img[ 5463] = 238;
assign img[ 5464] = 254;
assign img[ 5465] = 255;
assign img[ 5466] = 255;
assign img[ 5467] = 255;
assign img[ 5468] = 255;
assign img[ 5469] = 255;
assign img[ 5470] = 255;
assign img[ 5471] = 239;
assign img[ 5472] = 221;
assign img[ 5473] = 221;
assign img[ 5474] = 253;
assign img[ 5475] = 255;
assign img[ 5476] = 255;
assign img[ 5477] = 223;
assign img[ 5478] = 236;
assign img[ 5479] = 238;
assign img[ 5480] = 255;
assign img[ 5481] = 255;
assign img[ 5482] = 255;
assign img[ 5483] = 255;
assign img[ 5484] = 223;
assign img[ 5485] = 255;
assign img[ 5486] = 255;
assign img[ 5487] = 223;
assign img[ 5488] = 204;
assign img[ 5489] = 204;
assign img[ 5490] = 236;
assign img[ 5491] = 238;
assign img[ 5492] = 206;
assign img[ 5493] = 204;
assign img[ 5494] = 204;
assign img[ 5495] = 238;
assign img[ 5496] = 238;
assign img[ 5497] = 238;
assign img[ 5498] = 238;
assign img[ 5499] = 238;
assign img[ 5500] = 254;
assign img[ 5501] = 255;
assign img[ 5502] = 255;
assign img[ 5503] = 255;
assign img[ 5504] = 96;
assign img[ 5505] = 238;
assign img[ 5506] = 254;
assign img[ 5507] = 223;
assign img[ 5508] = 207;
assign img[ 5509] = 204;
assign img[ 5510] = 204;
assign img[ 5511] = 238;
assign img[ 5512] = 238;
assign img[ 5513] = 238;
assign img[ 5514] = 254;
assign img[ 5515] = 255;
assign img[ 5516] = 255;
assign img[ 5517] = 255;
assign img[ 5518] = 255;
assign img[ 5519] = 255;
assign img[ 5520] = 238;
assign img[ 5521] = 255;
assign img[ 5522] = 239;
assign img[ 5523] = 191;
assign img[ 5524] = 187;
assign img[ 5525] = 255;
assign img[ 5526] = 255;
assign img[ 5527] = 255;
assign img[ 5528] = 255;
assign img[ 5529] = 255;
assign img[ 5530] = 255;
assign img[ 5531] = 223;
assign img[ 5532] = 238;
assign img[ 5533] = 238;
assign img[ 5534] = 206;
assign img[ 5535] = 207;
assign img[ 5536] = 184;
assign img[ 5537] = 251;
assign img[ 5538] = 255;
assign img[ 5539] = 255;
assign img[ 5540] = 223;
assign img[ 5541] = 221;
assign img[ 5542] = 253;
assign img[ 5543] = 255;
assign img[ 5544] = 255;
assign img[ 5545] = 255;
assign img[ 5546] = 239;
assign img[ 5547] = 238;
assign img[ 5548] = 238;
assign img[ 5549] = 255;
assign img[ 5550] = 255;
assign img[ 5551] = 255;
assign img[ 5552] = 255;
assign img[ 5553] = 255;
assign img[ 5554] = 239;
assign img[ 5555] = 255;
assign img[ 5556] = 255;
assign img[ 5557] = 255;
assign img[ 5558] = 255;
assign img[ 5559] = 255;
assign img[ 5560] = 255;
assign img[ 5561] = 255;
assign img[ 5562] = 255;
assign img[ 5563] = 255;
assign img[ 5564] = 255;
assign img[ 5565] = 223;
assign img[ 5566] = 238;
assign img[ 5567] = 255;
assign img[ 5568] = 255;
assign img[ 5569] = 255;
assign img[ 5570] = 239;
assign img[ 5571] = 238;
assign img[ 5572] = 238;
assign img[ 5573] = 238;
assign img[ 5574] = 238;
assign img[ 5575] = 255;
assign img[ 5576] = 255;
assign img[ 5577] = 255;
assign img[ 5578] = 255;
assign img[ 5579] = 255;
assign img[ 5580] = 223;
assign img[ 5581] = 255;
assign img[ 5582] = 238;
assign img[ 5583] = 238;
assign img[ 5584] = 206;
assign img[ 5585] = 254;
assign img[ 5586] = 238;
assign img[ 5587] = 255;
assign img[ 5588] = 238;
assign img[ 5589] = 238;
assign img[ 5590] = 238;
assign img[ 5591] = 238;
assign img[ 5592] = 206;
assign img[ 5593] = 238;
assign img[ 5594] = 238;
assign img[ 5595] = 255;
assign img[ 5596] = 255;
assign img[ 5597] = 255;
assign img[ 5598] = 255;
assign img[ 5599] = 191;
assign img[ 5600] = 219;
assign img[ 5601] = 223;
assign img[ 5602] = 255;
assign img[ 5603] = 255;
assign img[ 5604] = 223;
assign img[ 5605] = 221;
assign img[ 5606] = 253;
assign img[ 5607] = 255;
assign img[ 5608] = 255;
assign img[ 5609] = 255;
assign img[ 5610] = 255;
assign img[ 5611] = 255;
assign img[ 5612] = 255;
assign img[ 5613] = 255;
assign img[ 5614] = 255;
assign img[ 5615] = 255;
assign img[ 5616] = 205;
assign img[ 5617] = 253;
assign img[ 5618] = 255;
assign img[ 5619] = 255;
assign img[ 5620] = 255;
assign img[ 5621] = 255;
assign img[ 5622] = 255;
assign img[ 5623] = 255;
assign img[ 5624] = 223;
assign img[ 5625] = 221;
assign img[ 5626] = 221;
assign img[ 5627] = 205;
assign img[ 5628] = 204;
assign img[ 5629] = 253;
assign img[ 5630] = 255;
assign img[ 5631] = 255;
assign img[ 5632] = 96;
assign img[ 5633] = 238;
assign img[ 5634] = 238;
assign img[ 5635] = 238;
assign img[ 5636] = 206;
assign img[ 5637] = 239;
assign img[ 5638] = 223;
assign img[ 5639] = 255;
assign img[ 5640] = 255;
assign img[ 5641] = 255;
assign img[ 5642] = 255;
assign img[ 5643] = 191;
assign img[ 5644] = 255;
assign img[ 5645] = 255;
assign img[ 5646] = 255;
assign img[ 5647] = 223;
assign img[ 5648] = 204;
assign img[ 5649] = 220;
assign img[ 5650] = 253;
assign img[ 5651] = 255;
assign img[ 5652] = 255;
assign img[ 5653] = 255;
assign img[ 5654] = 255;
assign img[ 5655] = 255;
assign img[ 5656] = 255;
assign img[ 5657] = 175;
assign img[ 5658] = 170;
assign img[ 5659] = 238;
assign img[ 5660] = 254;
assign img[ 5661] = 255;
assign img[ 5662] = 255;
assign img[ 5663] = 191;
assign img[ 5664] = 187;
assign img[ 5665] = 255;
assign img[ 5666] = 255;
assign img[ 5667] = 255;
assign img[ 5668] = 255;
assign img[ 5669] = 255;
assign img[ 5670] = 255;
assign img[ 5671] = 255;
assign img[ 5672] = 238;
assign img[ 5673] = 238;
assign img[ 5674] = 238;
assign img[ 5675] = 238;
assign img[ 5676] = 238;
assign img[ 5677] = 238;
assign img[ 5678] = 238;
assign img[ 5679] = 255;
assign img[ 5680] = 255;
assign img[ 5681] = 255;
assign img[ 5682] = 239;
assign img[ 5683] = 238;
assign img[ 5684] = 238;
assign img[ 5685] = 255;
assign img[ 5686] = 255;
assign img[ 5687] = 255;
assign img[ 5688] = 239;
assign img[ 5689] = 254;
assign img[ 5690] = 255;
assign img[ 5691] = 255;
assign img[ 5692] = 255;
assign img[ 5693] = 255;
assign img[ 5694] = 255;
assign img[ 5695] = 255;
assign img[ 5696] = 255;
assign img[ 5697] = 255;
assign img[ 5698] = 223;
assign img[ 5699] = 255;
assign img[ 5700] = 255;
assign img[ 5701] = 239;
assign img[ 5702] = 238;
assign img[ 5703] = 239;
assign img[ 5704] = 238;
assign img[ 5705] = 238;
assign img[ 5706] = 254;
assign img[ 5707] = 255;
assign img[ 5708] = 255;
assign img[ 5709] = 239;
assign img[ 5710] = 238;
assign img[ 5711] = 238;
assign img[ 5712] = 238;
assign img[ 5713] = 238;
assign img[ 5714] = 238;
assign img[ 5715] = 254;
assign img[ 5716] = 238;
assign img[ 5717] = 238;
assign img[ 5718] = 238;
assign img[ 5719] = 239;
assign img[ 5720] = 255;
assign img[ 5721] = 238;
assign img[ 5722] = 255;
assign img[ 5723] = 223;
assign img[ 5724] = 253;
assign img[ 5725] = 255;
assign img[ 5726] = 255;
assign img[ 5727] = 239;
assign img[ 5728] = 174;
assign img[ 5729] = 170;
assign img[ 5730] = 234;
assign img[ 5731] = 255;
assign img[ 5732] = 255;
assign img[ 5733] = 255;
assign img[ 5734] = 157;
assign img[ 5735] = 137;
assign img[ 5736] = 232;
assign img[ 5737] = 238;
assign img[ 5738] = 238;
assign img[ 5739] = 238;
assign img[ 5740] = 174;
assign img[ 5741] = 238;
assign img[ 5742] = 238;
assign img[ 5743] = 206;
assign img[ 5744] = 252;
assign img[ 5745] = 255;
assign img[ 5746] = 153;
assign img[ 5747] = 251;
assign img[ 5748] = 153;
assign img[ 5749] = 153;
assign img[ 5750] = 153;
assign img[ 5751] = 255;
assign img[ 5752] = 255;
assign img[ 5753] = 255;
assign img[ 5754] = 205;
assign img[ 5755] = 255;
assign img[ 5756] = 205;
assign img[ 5757] = 238;
assign img[ 5758] = 238;
assign img[ 5759] = 238;
assign img[ 5760] = 96;
assign img[ 5761] = 223;
assign img[ 5762] = 253;
assign img[ 5763] = 207;
assign img[ 5764] = 220;
assign img[ 5765] = 255;
assign img[ 5766] = 223;
assign img[ 5767] = 253;
assign img[ 5768] = 255;
assign img[ 5769] = 255;
assign img[ 5770] = 206;
assign img[ 5771] = 255;
assign img[ 5772] = 238;
assign img[ 5773] = 238;
assign img[ 5774] = 204;
assign img[ 5775] = 204;
assign img[ 5776] = 204;
assign img[ 5777] = 221;
assign img[ 5778] = 253;
assign img[ 5779] = 255;
assign img[ 5780] = 251;
assign img[ 5781] = 255;
assign img[ 5782] = 255;
assign img[ 5783] = 255;
assign img[ 5784] = 255;
assign img[ 5785] = 191;
assign img[ 5786] = 155;
assign img[ 5787] = 255;
assign img[ 5788] = 239;
assign img[ 5789] = 255;
assign img[ 5790] = 255;
assign img[ 5791] = 191;
assign img[ 5792] = 139;
assign img[ 5793] = 238;
assign img[ 5794] = 238;
assign img[ 5795] = 255;
assign img[ 5796] = 255;
assign img[ 5797] = 255;
assign img[ 5798] = 255;
assign img[ 5799] = 255;
assign img[ 5800] = 255;
assign img[ 5801] = 255;
assign img[ 5802] = 255;
assign img[ 5803] = 239;
assign img[ 5804] = 238;
assign img[ 5805] = 174;
assign img[ 5806] = 238;
assign img[ 5807] = 255;
assign img[ 5808] = 238;
assign img[ 5809] = 238;
assign img[ 5810] = 238;
assign img[ 5811] = 238;
assign img[ 5812] = 254;
assign img[ 5813] = 255;
assign img[ 5814] = 255;
assign img[ 5815] = 255;
assign img[ 5816] = 255;
assign img[ 5817] = 255;
assign img[ 5818] = 255;
assign img[ 5819] = 255;
assign img[ 5820] = 255;
assign img[ 5821] = 255;
assign img[ 5822] = 255;
assign img[ 5823] = 255;
assign img[ 5824] = 255;
assign img[ 5825] = 255;
assign img[ 5826] = 255;
assign img[ 5827] = 255;
assign img[ 5828] = 255;
assign img[ 5829] = 255;
assign img[ 5830] = 255;
assign img[ 5831] = 255;
assign img[ 5832] = 238;
assign img[ 5833] = 238;
assign img[ 5834] = 238;
assign img[ 5835] = 254;
assign img[ 5836] = 255;
assign img[ 5837] = 255;
assign img[ 5838] = 255;
assign img[ 5839] = 255;
assign img[ 5840] = 239;
assign img[ 5841] = 238;
assign img[ 5842] = 254;
assign img[ 5843] = 255;
assign img[ 5844] = 191;
assign img[ 5845] = 191;
assign img[ 5846] = 255;
assign img[ 5847] = 255;
assign img[ 5848] = 255;
assign img[ 5849] = 255;
assign img[ 5850] = 255;
assign img[ 5851] = 255;
assign img[ 5852] = 255;
assign img[ 5853] = 255;
assign img[ 5854] = 255;
assign img[ 5855] = 223;
assign img[ 5856] = 140;
assign img[ 5857] = 170;
assign img[ 5858] = 250;
assign img[ 5859] = 255;
assign img[ 5860] = 238;
assign img[ 5861] = 206;
assign img[ 5862] = 204;
assign img[ 5863] = 238;
assign img[ 5864] = 238;
assign img[ 5865] = 238;
assign img[ 5866] = 238;
assign img[ 5867] = 238;
assign img[ 5868] = 254;
assign img[ 5869] = 255;
assign img[ 5870] = 255;
assign img[ 5871] = 255;
assign img[ 5872] = 221;
assign img[ 5873] = 221;
assign img[ 5874] = 221;
assign img[ 5875] = 221;
assign img[ 5876] = 253;
assign img[ 5877] = 255;
assign img[ 5878] = 239;
assign img[ 5879] = 238;
assign img[ 5880] = 238;
assign img[ 5881] = 238;
assign img[ 5882] = 238;
assign img[ 5883] = 238;
assign img[ 5884] = 220;
assign img[ 5885] = 253;
assign img[ 5886] = 238;
assign img[ 5887] = 255;
assign img[ 5888] = 96;
assign img[ 5889] = 238;
assign img[ 5890] = 254;
assign img[ 5891] = 255;
assign img[ 5892] = 239;
assign img[ 5893] = 238;
assign img[ 5894] = 238;
assign img[ 5895] = 238;
assign img[ 5896] = 238;
assign img[ 5897] = 238;
assign img[ 5898] = 238;
assign img[ 5899] = 238;
assign img[ 5900] = 238;
assign img[ 5901] = 238;
assign img[ 5902] = 174;
assign img[ 5903] = 206;
assign img[ 5904] = 220;
assign img[ 5905] = 221;
assign img[ 5906] = 236;
assign img[ 5907] = 255;
assign img[ 5908] = 205;
assign img[ 5909] = 221;
assign img[ 5910] = 221;
assign img[ 5911] = 253;
assign img[ 5912] = 223;
assign img[ 5913] = 205;
assign img[ 5914] = 220;
assign img[ 5915] = 253;
assign img[ 5916] = 255;
assign img[ 5917] = 255;
assign img[ 5918] = 255;
assign img[ 5919] = 223;
assign img[ 5920] = 204;
assign img[ 5921] = 238;
assign img[ 5922] = 254;
assign img[ 5923] = 255;
assign img[ 5924] = 255;
assign img[ 5925] = 254;
assign img[ 5926] = 254;
assign img[ 5927] = 254;
assign img[ 5928] = 238;
assign img[ 5929] = 255;
assign img[ 5930] = 254;
assign img[ 5931] = 255;
assign img[ 5932] = 221;
assign img[ 5933] = 255;
assign img[ 5934] = 238;
assign img[ 5935] = 238;
assign img[ 5936] = 254;
assign img[ 5937] = 255;
assign img[ 5938] = 255;
assign img[ 5939] = 255;
assign img[ 5940] = 255;
assign img[ 5941] = 255;
assign img[ 5942] = 254;
assign img[ 5943] = 255;
assign img[ 5944] = 255;
assign img[ 5945] = 255;
assign img[ 5946] = 223;
assign img[ 5947] = 221;
assign img[ 5948] = 253;
assign img[ 5949] = 223;
assign img[ 5950] = 221;
assign img[ 5951] = 253;
assign img[ 5952] = 255;
assign img[ 5953] = 223;
assign img[ 5954] = 221;
assign img[ 5955] = 253;
assign img[ 5956] = 255;
assign img[ 5957] = 255;
assign img[ 5958] = 255;
assign img[ 5959] = 255;
assign img[ 5960] = 255;
assign img[ 5961] = 255;
assign img[ 5962] = 255;
assign img[ 5963] = 239;
assign img[ 5964] = 238;
assign img[ 5965] = 238;
assign img[ 5966] = 238;
assign img[ 5967] = 255;
assign img[ 5968] = 255;
assign img[ 5969] = 255;
assign img[ 5970] = 239;
assign img[ 5971] = 238;
assign img[ 5972] = 238;
assign img[ 5973] = 255;
assign img[ 5974] = 255;
assign img[ 5975] = 255;
assign img[ 5976] = 223;
assign img[ 5977] = 255;
assign img[ 5978] = 255;
assign img[ 5979] = 239;
assign img[ 5980] = 238;
assign img[ 5981] = 238;
assign img[ 5982] = 254;
assign img[ 5983] = 255;
assign img[ 5984] = 239;
assign img[ 5985] = 238;
assign img[ 5986] = 254;
assign img[ 5987] = 255;
assign img[ 5988] = 255;
assign img[ 5989] = 255;
assign img[ 5990] = 255;
assign img[ 5991] = 255;
assign img[ 5992] = 255;
assign img[ 5993] = 255;
assign img[ 5994] = 221;
assign img[ 5995] = 207;
assign img[ 5996] = 204;
assign img[ 5997] = 236;
assign img[ 5998] = 238;
assign img[ 5999] = 238;
assign img[ 6000] = 204;
assign img[ 6001] = 220;
assign img[ 6002] = 153;
assign img[ 6003] = 155;
assign img[ 6004] = 255;
assign img[ 6005] = 207;
assign img[ 6006] = 221;
assign img[ 6007] = 255;
assign img[ 6008] = 255;
assign img[ 6009] = 255;
assign img[ 6010] = 171;
assign img[ 6011] = 206;
assign img[ 6012] = 221;
assign img[ 6013] = 253;
assign img[ 6014] = 255;
assign img[ 6015] = 255;
assign img[ 6016] = 96;
assign img[ 6017] = 206;
assign img[ 6018] = 236;
assign img[ 6019] = 238;
assign img[ 6020] = 238;
assign img[ 6021] = 238;
assign img[ 6022] = 238;
assign img[ 6023] = 238;
assign img[ 6024] = 238;
assign img[ 6025] = 238;
assign img[ 6026] = 255;
assign img[ 6027] = 223;
assign img[ 6028] = 221;
assign img[ 6029] = 221;
assign img[ 6030] = 221;
assign img[ 6031] = 221;
assign img[ 6032] = 253;
assign img[ 6033] = 239;
assign img[ 6034] = 238;
assign img[ 6035] = 238;
assign img[ 6036] = 238;
assign img[ 6037] = 238;
assign img[ 6038] = 238;
assign img[ 6039] = 255;
assign img[ 6040] = 255;
assign img[ 6041] = 223;
assign img[ 6042] = 221;
assign img[ 6043] = 253;
assign img[ 6044] = 255;
assign img[ 6045] = 255;
assign img[ 6046] = 239;
assign img[ 6047] = 238;
assign img[ 6048] = 170;
assign img[ 6049] = 254;
assign img[ 6050] = 255;
assign img[ 6051] = 254;
assign img[ 6052] = 255;
assign img[ 6053] = 255;
assign img[ 6054] = 255;
assign img[ 6055] = 255;
assign img[ 6056] = 238;
assign img[ 6057] = 238;
assign img[ 6058] = 254;
assign img[ 6059] = 191;
assign img[ 6060] = 187;
assign img[ 6061] = 255;
assign img[ 6062] = 238;
assign img[ 6063] = 255;
assign img[ 6064] = 255;
assign img[ 6065] = 255;
assign img[ 6066] = 255;
assign img[ 6067] = 255;
assign img[ 6068] = 255;
assign img[ 6069] = 255;
assign img[ 6070] = 255;
assign img[ 6071] = 255;
assign img[ 6072] = 223;
assign img[ 6073] = 221;
assign img[ 6074] = 221;
assign img[ 6075] = 255;
assign img[ 6076] = 255;
assign img[ 6077] = 207;
assign img[ 6078] = 238;
assign img[ 6079] = 255;
assign img[ 6080] = 255;
assign img[ 6081] = 255;
assign img[ 6082] = 223;
assign img[ 6083] = 255;
assign img[ 6084] = 255;
assign img[ 6085] = 255;
assign img[ 6086] = 255;
assign img[ 6087] = 223;
assign img[ 6088] = 253;
assign img[ 6089] = 255;
assign img[ 6090] = 255;
assign img[ 6091] = 239;
assign img[ 6092] = 238;
assign img[ 6093] = 238;
assign img[ 6094] = 238;
assign img[ 6095] = 255;
assign img[ 6096] = 255;
assign img[ 6097] = 255;
assign img[ 6098] = 239;
assign img[ 6099] = 254;
assign img[ 6100] = 191;
assign img[ 6101] = 255;
assign img[ 6102] = 255;
assign img[ 6103] = 255;
assign img[ 6104] = 239;
assign img[ 6105] = 238;
assign img[ 6106] = 238;
assign img[ 6107] = 238;
assign img[ 6108] = 238;
assign img[ 6109] = 238;
assign img[ 6110] = 255;
assign img[ 6111] = 255;
assign img[ 6112] = 255;
assign img[ 6113] = 255;
assign img[ 6114] = 238;
assign img[ 6115] = 238;
assign img[ 6116] = 238;
assign img[ 6117] = 238;
assign img[ 6118] = 238;
assign img[ 6119] = 238;
assign img[ 6120] = 254;
assign img[ 6121] = 255;
assign img[ 6122] = 255;
assign img[ 6123] = 255;
assign img[ 6124] = 255;
assign img[ 6125] = 255;
assign img[ 6126] = 255;
assign img[ 6127] = 255;
assign img[ 6128] = 223;
assign img[ 6129] = 221;
assign img[ 6130] = 185;
assign img[ 6131] = 255;
assign img[ 6132] = 223;
assign img[ 6133] = 221;
assign img[ 6134] = 253;
assign img[ 6135] = 255;
assign img[ 6136] = 255;
assign img[ 6137] = 207;
assign img[ 6138] = 204;
assign img[ 6139] = 221;
assign img[ 6140] = 253;
assign img[ 6141] = 255;
assign img[ 6142] = 255;
assign img[ 6143] = 255;
assign img[ 6144] = 96;
assign img[ 6145] = 255;
assign img[ 6146] = 255;
assign img[ 6147] = 223;
assign img[ 6148] = 205;
assign img[ 6149] = 238;
assign img[ 6150] = 238;
assign img[ 6151] = 238;
assign img[ 6152] = 238;
assign img[ 6153] = 238;
assign img[ 6154] = 254;
assign img[ 6155] = 175;
assign img[ 6156] = 170;
assign img[ 6157] = 238;
assign img[ 6158] = 238;
assign img[ 6159] = 239;
assign img[ 6160] = 238;
assign img[ 6161] = 238;
assign img[ 6162] = 238;
assign img[ 6163] = 174;
assign img[ 6164] = 170;
assign img[ 6165] = 238;
assign img[ 6166] = 238;
assign img[ 6167] = 238;
assign img[ 6168] = 238;
assign img[ 6169] = 238;
assign img[ 6170] = 204;
assign img[ 6171] = 238;
assign img[ 6172] = 238;
assign img[ 6173] = 255;
assign img[ 6174] = 223;
assign img[ 6175] = 159;
assign img[ 6176] = 185;
assign img[ 6177] = 238;
assign img[ 6178] = 222;
assign img[ 6179] = 253;
assign img[ 6180] = 255;
assign img[ 6181] = 255;
assign img[ 6182] = 255;
assign img[ 6183] = 255;
assign img[ 6184] = 238;
assign img[ 6185] = 238;
assign img[ 6186] = 255;
assign img[ 6187] = 254;
assign img[ 6188] = 238;
assign img[ 6189] = 223;
assign img[ 6190] = 254;
assign img[ 6191] = 255;
assign img[ 6192] = 255;
assign img[ 6193] = 255;
assign img[ 6194] = 255;
assign img[ 6195] = 255;
assign img[ 6196] = 255;
assign img[ 6197] = 255;
assign img[ 6198] = 255;
assign img[ 6199] = 255;
assign img[ 6200] = 255;
assign img[ 6201] = 223;
assign img[ 6202] = 238;
assign img[ 6203] = 238;
assign img[ 6204] = 238;
assign img[ 6205] = 255;
assign img[ 6206] = 255;
assign img[ 6207] = 255;
assign img[ 6208] = 255;
assign img[ 6209] = 255;
assign img[ 6210] = 255;
assign img[ 6211] = 255;
assign img[ 6212] = 255;
assign img[ 6213] = 255;
assign img[ 6214] = 139;
assign img[ 6215] = 238;
assign img[ 6216] = 254;
assign img[ 6217] = 255;
assign img[ 6218] = 255;
assign img[ 6219] = 255;
assign img[ 6220] = 255;
assign img[ 6221] = 239;
assign img[ 6222] = 204;
assign img[ 6223] = 254;
assign img[ 6224] = 255;
assign img[ 6225] = 255;
assign img[ 6226] = 255;
assign img[ 6227] = 255;
assign img[ 6228] = 255;
assign img[ 6229] = 207;
assign img[ 6230] = 238;
assign img[ 6231] = 238;
assign img[ 6232] = 238;
assign img[ 6233] = 238;
assign img[ 6234] = 254;
assign img[ 6235] = 255;
assign img[ 6236] = 255;
assign img[ 6237] = 255;
assign img[ 6238] = 238;
assign img[ 6239] = 206;
assign img[ 6240] = 156;
assign img[ 6241] = 153;
assign img[ 6242] = 249;
assign img[ 6243] = 255;
assign img[ 6244] = 255;
assign img[ 6245] = 255;
assign img[ 6246] = 223;
assign img[ 6247] = 255;
assign img[ 6248] = 255;
assign img[ 6249] = 255;
assign img[ 6250] = 238;
assign img[ 6251] = 255;
assign img[ 6252] = 255;
assign img[ 6253] = 255;
assign img[ 6254] = 255;
assign img[ 6255] = 255;
assign img[ 6256] = 171;
assign img[ 6257] = 238;
assign img[ 6258] = 238;
assign img[ 6259] = 255;
assign img[ 6260] = 191;
assign img[ 6261] = 155;
assign img[ 6262] = 217;
assign img[ 6263] = 255;
assign img[ 6264] = 255;
assign img[ 6265] = 255;
assign img[ 6266] = 238;
assign img[ 6267] = 238;
assign img[ 6268] = 254;
assign img[ 6269] = 255;
assign img[ 6270] = 223;
assign img[ 6271] = 255;
assign img[ 6272] = 96;
assign img[ 6273] = 206;
assign img[ 6274] = 236;
assign img[ 6275] = 223;
assign img[ 6276] = 205;
assign img[ 6277] = 236;
assign img[ 6278] = 206;
assign img[ 6279] = 236;
assign img[ 6280] = 238;
assign img[ 6281] = 238;
assign img[ 6282] = 238;
assign img[ 6283] = 206;
assign img[ 6284] = 204;
assign img[ 6285] = 221;
assign img[ 6286] = 221;
assign img[ 6287] = 221;
assign img[ 6288] = 204;
assign img[ 6289] = 204;
assign img[ 6290] = 236;
assign img[ 6291] = 238;
assign img[ 6292] = 238;
assign img[ 6293] = 254;
assign img[ 6294] = 206;
assign img[ 6295] = 252;
assign img[ 6296] = 254;
assign img[ 6297] = 255;
assign img[ 6298] = 187;
assign img[ 6299] = 255;
assign img[ 6300] = 223;
assign img[ 6301] = 255;
assign img[ 6302] = 255;
assign img[ 6303] = 255;
assign img[ 6304] = 155;
assign img[ 6305] = 169;
assign img[ 6306] = 238;
assign img[ 6307] = 238;
assign img[ 6308] = 238;
assign img[ 6309] = 238;
assign img[ 6310] = 238;
assign img[ 6311] = 238;
assign img[ 6312] = 238;
assign img[ 6313] = 238;
assign img[ 6314] = 238;
assign img[ 6315] = 238;
assign img[ 6316] = 238;
assign img[ 6317] = 222;
assign img[ 6318] = 253;
assign img[ 6319] = 238;
assign img[ 6320] = 238;
assign img[ 6321] = 238;
assign img[ 6322] = 204;
assign img[ 6323] = 238;
assign img[ 6324] = 238;
assign img[ 6325] = 238;
assign img[ 6326] = 238;
assign img[ 6327] = 238;
assign img[ 6328] = 238;
assign img[ 6329] = 238;
assign img[ 6330] = 238;
assign img[ 6331] = 238;
assign img[ 6332] = 238;
assign img[ 6333] = 254;
assign img[ 6334] = 255;
assign img[ 6335] = 255;
assign img[ 6336] = 238;
assign img[ 6337] = 254;
assign img[ 6338] = 238;
assign img[ 6339] = 238;
assign img[ 6340] = 206;
assign img[ 6341] = 204;
assign img[ 6342] = 204;
assign img[ 6343] = 204;
assign img[ 6344] = 236;
assign img[ 6345] = 238;
assign img[ 6346] = 238;
assign img[ 6347] = 255;
assign img[ 6348] = 238;
assign img[ 6349] = 239;
assign img[ 6350] = 255;
assign img[ 6351] = 254;
assign img[ 6352] = 255;
assign img[ 6353] = 255;
assign img[ 6354] = 254;
assign img[ 6355] = 255;
assign img[ 6356] = 238;
assign img[ 6357] = 207;
assign img[ 6358] = 238;
assign img[ 6359] = 238;
assign img[ 6360] = 238;
assign img[ 6361] = 238;
assign img[ 6362] = 238;
assign img[ 6363] = 238;
assign img[ 6364] = 254;
assign img[ 6365] = 255;
assign img[ 6366] = 239;
assign img[ 6367] = 206;
assign img[ 6368] = 204;
assign img[ 6369] = 221;
assign img[ 6370] = 253;
assign img[ 6371] = 255;
assign img[ 6372] = 255;
assign img[ 6373] = 255;
assign img[ 6374] = 255;
assign img[ 6375] = 255;
assign img[ 6376] = 255;
assign img[ 6377] = 255;
assign img[ 6378] = 255;
assign img[ 6379] = 255;
assign img[ 6380] = 255;
assign img[ 6381] = 255;
assign img[ 6382] = 255;
assign img[ 6383] = 255;
assign img[ 6384] = 239;
assign img[ 6385] = 206;
assign img[ 6386] = 220;
assign img[ 6387] = 223;
assign img[ 6388] = 253;
assign img[ 6389] = 255;
assign img[ 6390] = 238;
assign img[ 6391] = 238;
assign img[ 6392] = 238;
assign img[ 6393] = 238;
assign img[ 6394] = 238;
assign img[ 6395] = 207;
assign img[ 6396] = 236;
assign img[ 6397] = 238;
assign img[ 6398] = 222;
assign img[ 6399] = 255;
assign img[ 6400] = 96;
assign img[ 6401] = 238;
assign img[ 6402] = 238;
assign img[ 6403] = 255;
assign img[ 6404] = 239;
assign img[ 6405] = 255;
assign img[ 6406] = 239;
assign img[ 6407] = 238;
assign img[ 6408] = 238;
assign img[ 6409] = 238;
assign img[ 6410] = 238;
assign img[ 6411] = 223;
assign img[ 6412] = 221;
assign img[ 6413] = 253;
assign img[ 6414] = 255;
assign img[ 6415] = 223;
assign img[ 6416] = 221;
assign img[ 6417] = 205;
assign img[ 6418] = 236;
assign img[ 6419] = 239;
assign img[ 6420] = 204;
assign img[ 6421] = 238;
assign img[ 6422] = 238;
assign img[ 6423] = 238;
assign img[ 6424] = 238;
assign img[ 6425] = 254;
assign img[ 6426] = 187;
assign img[ 6427] = 255;
assign img[ 6428] = 255;
assign img[ 6429] = 255;
assign img[ 6430] = 239;
assign img[ 6431] = 174;
assign img[ 6432] = 186;
assign img[ 6433] = 255;
assign img[ 6434] = 255;
assign img[ 6435] = 255;
assign img[ 6436] = 255;
assign img[ 6437] = 255;
assign img[ 6438] = 255;
assign img[ 6439] = 239;
assign img[ 6440] = 238;
assign img[ 6441] = 238;
assign img[ 6442] = 238;
assign img[ 6443] = 238;
assign img[ 6444] = 238;
assign img[ 6445] = 254;
assign img[ 6446] = 255;
assign img[ 6447] = 255;
assign img[ 6448] = 255;
assign img[ 6449] = 255;
assign img[ 6450] = 239;
assign img[ 6451] = 238;
assign img[ 6452] = 238;
assign img[ 6453] = 255;
assign img[ 6454] = 255;
assign img[ 6455] = 239;
assign img[ 6456] = 238;
assign img[ 6457] = 238;
assign img[ 6458] = 254;
assign img[ 6459] = 255;
assign img[ 6460] = 255;
assign img[ 6461] = 255;
assign img[ 6462] = 255;
assign img[ 6463] = 255;
assign img[ 6464] = 255;
assign img[ 6465] = 255;
assign img[ 6466] = 255;
assign img[ 6467] = 255;
assign img[ 6468] = 255;
assign img[ 6469] = 255;
assign img[ 6470] = 255;
assign img[ 6471] = 255;
assign img[ 6472] = 255;
assign img[ 6473] = 255;
assign img[ 6474] = 255;
assign img[ 6475] = 255;
assign img[ 6476] = 255;
assign img[ 6477] = 255;
assign img[ 6478] = 238;
assign img[ 6479] = 255;
assign img[ 6480] = 255;
assign img[ 6481] = 255;
assign img[ 6482] = 255;
assign img[ 6483] = 255;
assign img[ 6484] = 238;
assign img[ 6485] = 238;
assign img[ 6486] = 238;
assign img[ 6487] = 238;
assign img[ 6488] = 238;
assign img[ 6489] = 238;
assign img[ 6490] = 238;
assign img[ 6491] = 255;
assign img[ 6492] = 255;
assign img[ 6493] = 255;
assign img[ 6494] = 255;
assign img[ 6495] = 255;
assign img[ 6496] = 171;
assign img[ 6497] = 170;
assign img[ 6498] = 250;
assign img[ 6499] = 255;
assign img[ 6500] = 255;
assign img[ 6501] = 255;
assign img[ 6502] = 255;
assign img[ 6503] = 255;
assign img[ 6504] = 239;
assign img[ 6505] = 238;
assign img[ 6506] = 238;
assign img[ 6507] = 238;
assign img[ 6508] = 206;
assign img[ 6509] = 238;
assign img[ 6510] = 238;
assign img[ 6511] = 206;
assign img[ 6512] = 204;
assign img[ 6513] = 236;
assign img[ 6514] = 238;
assign img[ 6515] = 255;
assign img[ 6516] = 207;
assign img[ 6517] = 223;
assign img[ 6518] = 255;
assign img[ 6519] = 255;
assign img[ 6520] = 255;
assign img[ 6521] = 239;
assign img[ 6522] = 254;
assign img[ 6523] = 239;
assign img[ 6524] = 238;
assign img[ 6525] = 238;
assign img[ 6526] = 238;
assign img[ 6527] = 238;
assign img[ 6528] = 0;
assign img[ 6529] = 186;
assign img[ 6530] = 251;
assign img[ 6531] = 255;
assign img[ 6532] = 255;
assign img[ 6533] = 255;
assign img[ 6534] = 255;
assign img[ 6535] = 255;
assign img[ 6536] = 255;
assign img[ 6537] = 255;
assign img[ 6538] = 255;
assign img[ 6539] = 239;
assign img[ 6540] = 238;
assign img[ 6541] = 238;
assign img[ 6542] = 254;
assign img[ 6543] = 239;
assign img[ 6544] = 206;
assign img[ 6545] = 238;
assign img[ 6546] = 254;
assign img[ 6547] = 255;
assign img[ 6548] = 255;
assign img[ 6549] = 255;
assign img[ 6550] = 238;
assign img[ 6551] = 254;
assign img[ 6552] = 255;
assign img[ 6553] = 238;
assign img[ 6554] = 204;
assign img[ 6555] = 204;
assign img[ 6556] = 236;
assign img[ 6557] = 238;
assign img[ 6558] = 223;
assign img[ 6559] = 205;
assign img[ 6560] = 204;
assign img[ 6561] = 255;
assign img[ 6562] = 255;
assign img[ 6563] = 255;
assign img[ 6564] = 255;
assign img[ 6565] = 255;
assign img[ 6566] = 255;
assign img[ 6567] = 255;
assign img[ 6568] = 238;
assign img[ 6569] = 238;
assign img[ 6570] = 255;
assign img[ 6571] = 255;
assign img[ 6572] = 255;
assign img[ 6573] = 223;
assign img[ 6574] = 253;
assign img[ 6575] = 239;
assign img[ 6576] = 238;
assign img[ 6577] = 239;
assign img[ 6578] = 238;
assign img[ 6579] = 238;
assign img[ 6580] = 238;
assign img[ 6581] = 238;
assign img[ 6582] = 238;
assign img[ 6583] = 238;
assign img[ 6584] = 238;
assign img[ 6585] = 254;
assign img[ 6586] = 254;
assign img[ 6587] = 255;
assign img[ 6588] = 255;
assign img[ 6589] = 255;
assign img[ 6590] = 239;
assign img[ 6591] = 238;
assign img[ 6592] = 238;
assign img[ 6593] = 207;
assign img[ 6594] = 220;
assign img[ 6595] = 255;
assign img[ 6596] = 255;
assign img[ 6597] = 255;
assign img[ 6598] = 255;
assign img[ 6599] = 255;
assign img[ 6600] = 255;
assign img[ 6601] = 255;
assign img[ 6602] = 255;
assign img[ 6603] = 255;
assign img[ 6604] = 255;
assign img[ 6605] = 255;
assign img[ 6606] = 239;
assign img[ 6607] = 238;
assign img[ 6608] = 206;
assign img[ 6609] = 238;
assign img[ 6610] = 254;
assign img[ 6611] = 255;
assign img[ 6612] = 239;
assign img[ 6613] = 238;
assign img[ 6614] = 238;
assign img[ 6615] = 238;
assign img[ 6616] = 238;
assign img[ 6617] = 238;
assign img[ 6618] = 238;
assign img[ 6619] = 255;
assign img[ 6620] = 238;
assign img[ 6621] = 255;
assign img[ 6622] = 255;
assign img[ 6623] = 255;
assign img[ 6624] = 187;
assign img[ 6625] = 255;
assign img[ 6626] = 255;
assign img[ 6627] = 255;
assign img[ 6628] = 255;
assign img[ 6629] = 255;
assign img[ 6630] = 255;
assign img[ 6631] = 255;
assign img[ 6632] = 255;
assign img[ 6633] = 255;
assign img[ 6634] = 238;
assign img[ 6635] = 238;
assign img[ 6636] = 238;
assign img[ 6637] = 238;
assign img[ 6638] = 238;
assign img[ 6639] = 255;
assign img[ 6640] = 221;
assign img[ 6641] = 255;
assign img[ 6642] = 255;
assign img[ 6643] = 239;
assign img[ 6644] = 206;
assign img[ 6645] = 204;
assign img[ 6646] = 204;
assign img[ 6647] = 238;
assign img[ 6648] = 238;
assign img[ 6649] = 206;
assign img[ 6650] = 204;
assign img[ 6651] = 221;
assign img[ 6652] = 205;
assign img[ 6653] = 238;
assign img[ 6654] = 206;
assign img[ 6655] = 204;
assign img[ 6656] = 96;
assign img[ 6657] = 239;
assign img[ 6658] = 238;
assign img[ 6659] = 238;
assign img[ 6660] = 206;
assign img[ 6661] = 220;
assign img[ 6662] = 221;
assign img[ 6663] = 253;
assign img[ 6664] = 255;
assign img[ 6665] = 255;
assign img[ 6666] = 255;
assign img[ 6667] = 255;
assign img[ 6668] = 255;
assign img[ 6669] = 239;
assign img[ 6670] = 238;
assign img[ 6671] = 255;
assign img[ 6672] = 255;
assign img[ 6673] = 255;
assign img[ 6674] = 238;
assign img[ 6675] = 255;
assign img[ 6676] = 239;
assign img[ 6677] = 238;
assign img[ 6678] = 206;
assign img[ 6679] = 238;
assign img[ 6680] = 238;
assign img[ 6681] = 191;
assign img[ 6682] = 187;
assign img[ 6683] = 251;
assign img[ 6684] = 255;
assign img[ 6685] = 255;
assign img[ 6686] = 254;
assign img[ 6687] = 255;
assign img[ 6688] = 255;
assign img[ 6689] = 255;
assign img[ 6690] = 239;
assign img[ 6691] = 238;
assign img[ 6692] = 238;
assign img[ 6693] = 238;
assign img[ 6694] = 238;
assign img[ 6695] = 255;
assign img[ 6696] = 255;
assign img[ 6697] = 255;
assign img[ 6698] = 239;
assign img[ 6699] = 238;
assign img[ 6700] = 238;
assign img[ 6701] = 254;
assign img[ 6702] = 255;
assign img[ 6703] = 238;
assign img[ 6704] = 254;
assign img[ 6705] = 255;
assign img[ 6706] = 255;
assign img[ 6707] = 255;
assign img[ 6708] = 238;
assign img[ 6709] = 255;
assign img[ 6710] = 254;
assign img[ 6711] = 255;
assign img[ 6712] = 254;
assign img[ 6713] = 255;
assign img[ 6714] = 255;
assign img[ 6715] = 255;
assign img[ 6716] = 255;
assign img[ 6717] = 223;
assign img[ 6718] = 255;
assign img[ 6719] = 255;
assign img[ 6720] = 255;
assign img[ 6721] = 255;
assign img[ 6722] = 255;
assign img[ 6723] = 255;
assign img[ 6724] = 255;
assign img[ 6725] = 255;
assign img[ 6726] = 255;
assign img[ 6727] = 255;
assign img[ 6728] = 255;
assign img[ 6729] = 255;
assign img[ 6730] = 255;
assign img[ 6731] = 255;
assign img[ 6732] = 255;
assign img[ 6733] = 255;
assign img[ 6734] = 255;
assign img[ 6735] = 255;
assign img[ 6736] = 255;
assign img[ 6737] = 255;
assign img[ 6738] = 255;
assign img[ 6739] = 239;
assign img[ 6740] = 238;
assign img[ 6741] = 239;
assign img[ 6742] = 238;
assign img[ 6743] = 238;
assign img[ 6744] = 238;
assign img[ 6745] = 238;
assign img[ 6746] = 238;
assign img[ 6747] = 255;
assign img[ 6748] = 238;
assign img[ 6749] = 239;
assign img[ 6750] = 238;
assign img[ 6751] = 238;
assign img[ 6752] = 220;
assign img[ 6753] = 253;
assign img[ 6754] = 238;
assign img[ 6755] = 238;
assign img[ 6756] = 238;
assign img[ 6757] = 191;
assign img[ 6758] = 187;
assign img[ 6759] = 251;
assign img[ 6760] = 255;
assign img[ 6761] = 255;
assign img[ 6762] = 238;
assign img[ 6763] = 238;
assign img[ 6764] = 238;
assign img[ 6765] = 238;
assign img[ 6766] = 238;
assign img[ 6767] = 238;
assign img[ 6768] = 238;
assign img[ 6769] = 238;
assign img[ 6770] = 238;
assign img[ 6771] = 222;
assign img[ 6772] = 205;
assign img[ 6773] = 223;
assign img[ 6774] = 255;
assign img[ 6775] = 239;
assign img[ 6776] = 238;
assign img[ 6777] = 238;
assign img[ 6778] = 238;
assign img[ 6779] = 223;
assign img[ 6780] = 253;
assign img[ 6781] = 254;
assign img[ 6782] = 238;
assign img[ 6783] = 238;
assign img[ 6784] = 96;
assign img[ 6785] = 255;
assign img[ 6786] = 255;
assign img[ 6787] = 255;
assign img[ 6788] = 255;
assign img[ 6789] = 255;
assign img[ 6790] = 255;
assign img[ 6791] = 255;
assign img[ 6792] = 238;
assign img[ 6793] = 254;
assign img[ 6794] = 254;
assign img[ 6795] = 223;
assign img[ 6796] = 204;
assign img[ 6797] = 236;
assign img[ 6798] = 206;
assign img[ 6799] = 205;
assign img[ 6800] = 221;
assign img[ 6801] = 255;
assign img[ 6802] = 255;
assign img[ 6803] = 255;
assign img[ 6804] = 255;
assign img[ 6805] = 255;
assign img[ 6806] = 255;
assign img[ 6807] = 255;
assign img[ 6808] = 255;
assign img[ 6809] = 255;
assign img[ 6810] = 255;
assign img[ 6811] = 255;
assign img[ 6812] = 255;
assign img[ 6813] = 255;
assign img[ 6814] = 239;
assign img[ 6815] = 255;
assign img[ 6816] = 255;
assign img[ 6817] = 255;
assign img[ 6818] = 255;
assign img[ 6819] = 255;
assign img[ 6820] = 239;
assign img[ 6821] = 239;
assign img[ 6822] = 255;
assign img[ 6823] = 255;
assign img[ 6824] = 255;
assign img[ 6825] = 255;
assign img[ 6826] = 255;
assign img[ 6827] = 255;
assign img[ 6828] = 223;
assign img[ 6829] = 223;
assign img[ 6830] = 238;
assign img[ 6831] = 255;
assign img[ 6832] = 255;
assign img[ 6833] = 255;
assign img[ 6834] = 255;
assign img[ 6835] = 255;
assign img[ 6836] = 255;
assign img[ 6837] = 255;
assign img[ 6838] = 239;
assign img[ 6839] = 238;
assign img[ 6840] = 238;
assign img[ 6841] = 238;
assign img[ 6842] = 238;
assign img[ 6843] = 254;
assign img[ 6844] = 255;
assign img[ 6845] = 255;
assign img[ 6846] = 238;
assign img[ 6847] = 255;
assign img[ 6848] = 255;
assign img[ 6849] = 255;
assign img[ 6850] = 239;
assign img[ 6851] = 255;
assign img[ 6852] = 255;
assign img[ 6853] = 239;
assign img[ 6854] = 238;
assign img[ 6855] = 238;
assign img[ 6856] = 238;
assign img[ 6857] = 238;
assign img[ 6858] = 254;
assign img[ 6859] = 255;
assign img[ 6860] = 255;
assign img[ 6861] = 239;
assign img[ 6862] = 238;
assign img[ 6863] = 255;
assign img[ 6864] = 255;
assign img[ 6865] = 255;
assign img[ 6866] = 239;
assign img[ 6867] = 222;
assign img[ 6868] = 253;
assign img[ 6869] = 255;
assign img[ 6870] = 255;
assign img[ 6871] = 223;
assign img[ 6872] = 221;
assign img[ 6873] = 253;
assign img[ 6874] = 255;
assign img[ 6875] = 255;
assign img[ 6876] = 255;
assign img[ 6877] = 255;
assign img[ 6878] = 255;
assign img[ 6879] = 255;
assign img[ 6880] = 221;
assign img[ 6881] = 221;
assign img[ 6882] = 253;
assign img[ 6883] = 255;
assign img[ 6884] = 255;
assign img[ 6885] = 223;
assign img[ 6886] = 221;
assign img[ 6887] = 255;
assign img[ 6888] = 255;
assign img[ 6889] = 255;
assign img[ 6890] = 255;
assign img[ 6891] = 239;
assign img[ 6892] = 238;
assign img[ 6893] = 238;
assign img[ 6894] = 238;
assign img[ 6895] = 238;
assign img[ 6896] = 238;
assign img[ 6897] = 206;
assign img[ 6898] = 236;
assign img[ 6899] = 239;
assign img[ 6900] = 204;
assign img[ 6901] = 236;
assign img[ 6902] = 238;
assign img[ 6903] = 238;
assign img[ 6904] = 238;
assign img[ 6905] = 174;
assign img[ 6906] = 170;
assign img[ 6907] = 238;
assign img[ 6908] = 238;
assign img[ 6909] = 255;
assign img[ 6910] = 255;
assign img[ 6911] = 255;
assign img[ 6912] = 96;
assign img[ 6913] = 238;
assign img[ 6914] = 238;
assign img[ 6915] = 238;
assign img[ 6916] = 255;
assign img[ 6917] = 255;
assign img[ 6918] = 239;
assign img[ 6919] = 238;
assign img[ 6920] = 238;
assign img[ 6921] = 238;
assign img[ 6922] = 238;
assign img[ 6923] = 206;
assign img[ 6924] = 204;
assign img[ 6925] = 204;
assign img[ 6926] = 220;
assign img[ 6927] = 221;
assign img[ 6928] = 221;
assign img[ 6929] = 253;
assign img[ 6930] = 255;
assign img[ 6931] = 191;
assign img[ 6932] = 171;
assign img[ 6933] = 238;
assign img[ 6934] = 238;
assign img[ 6935] = 238;
assign img[ 6936] = 238;
assign img[ 6937] = 223;
assign img[ 6938] = 221;
assign img[ 6939] = 221;
assign img[ 6940] = 253;
assign img[ 6941] = 255;
assign img[ 6942] = 255;
assign img[ 6943] = 255;
assign img[ 6944] = 187;
assign img[ 6945] = 251;
assign img[ 6946] = 255;
assign img[ 6947] = 255;
assign img[ 6948] = 255;
assign img[ 6949] = 239;
assign img[ 6950] = 238;
assign img[ 6951] = 239;
assign img[ 6952] = 238;
assign img[ 6953] = 238;
assign img[ 6954] = 206;
assign img[ 6955] = 238;
assign img[ 6956] = 238;
assign img[ 6957] = 238;
assign img[ 6958] = 238;
assign img[ 6959] = 238;
assign img[ 6960] = 254;
assign img[ 6961] = 255;
assign img[ 6962] = 255;
assign img[ 6963] = 207;
assign img[ 6964] = 236;
assign img[ 6965] = 255;
assign img[ 6966] = 255;
assign img[ 6967] = 255;
assign img[ 6968] = 239;
assign img[ 6969] = 238;
assign img[ 6970] = 254;
assign img[ 6971] = 255;
assign img[ 6972] = 255;
assign img[ 6973] = 239;
assign img[ 6974] = 238;
assign img[ 6975] = 255;
assign img[ 6976] = 255;
assign img[ 6977] = 255;
assign img[ 6978] = 223;
assign img[ 6979] = 255;
assign img[ 6980] = 255;
assign img[ 6981] = 255;
assign img[ 6982] = 255;
assign img[ 6983] = 255;
assign img[ 6984] = 238;
assign img[ 6985] = 238;
assign img[ 6986] = 254;
assign img[ 6987] = 255;
assign img[ 6988] = 255;
assign img[ 6989] = 255;
assign img[ 6990] = 255;
assign img[ 6991] = 255;
assign img[ 6992] = 255;
assign img[ 6993] = 255;
assign img[ 6994] = 255;
assign img[ 6995] = 255;
assign img[ 6996] = 255;
assign img[ 6997] = 255;
assign img[ 6998] = 238;
assign img[ 6999] = 238;
assign img[ 7000] = 255;
assign img[ 7001] = 255;
assign img[ 7002] = 206;
assign img[ 7003] = 238;
assign img[ 7004] = 254;
assign img[ 7005] = 255;
assign img[ 7006] = 255;
assign img[ 7007] = 191;
assign img[ 7008] = 234;
assign img[ 7009] = 255;
assign img[ 7010] = 255;
assign img[ 7011] = 255;
assign img[ 7012] = 223;
assign img[ 7013] = 221;
assign img[ 7014] = 221;
assign img[ 7015] = 221;
assign img[ 7016] = 253;
assign img[ 7017] = 255;
assign img[ 7018] = 255;
assign img[ 7019] = 239;
assign img[ 7020] = 204;
assign img[ 7021] = 238;
assign img[ 7022] = 238;
assign img[ 7023] = 238;
assign img[ 7024] = 254;
assign img[ 7025] = 255;
assign img[ 7026] = 221;
assign img[ 7027] = 191;
assign img[ 7028] = 139;
assign img[ 7029] = 204;
assign img[ 7030] = 236;
assign img[ 7031] = 238;
assign img[ 7032] = 238;
assign img[ 7033] = 174;
assign img[ 7034] = 238;
assign img[ 7035] = 238;
assign img[ 7036] = 220;
assign img[ 7037] = 253;
assign img[ 7038] = 255;
assign img[ 7039] = 255;
assign img[ 7040] = 96;
assign img[ 7041] = 191;
assign img[ 7042] = 251;
assign img[ 7043] = 255;
assign img[ 7044] = 187;
assign img[ 7045] = 187;
assign img[ 7046] = 187;
assign img[ 7047] = 251;
assign img[ 7048] = 255;
assign img[ 7049] = 255;
assign img[ 7050] = 239;
assign img[ 7051] = 190;
assign img[ 7052] = 255;
assign img[ 7053] = 255;
assign img[ 7054] = 255;
assign img[ 7055] = 255;
assign img[ 7056] = 238;
assign img[ 7057] = 223;
assign img[ 7058] = 221;
assign img[ 7059] = 223;
assign img[ 7060] = 221;
assign img[ 7061] = 255;
assign img[ 7062] = 223;
assign img[ 7063] = 253;
assign img[ 7064] = 254;
assign img[ 7065] = 174;
assign img[ 7066] = 186;
assign img[ 7067] = 255;
assign img[ 7068] = 255;
assign img[ 7069] = 255;
assign img[ 7070] = 238;
assign img[ 7071] = 206;
assign img[ 7072] = 204;
assign img[ 7073] = 253;
assign img[ 7074] = 255;
assign img[ 7075] = 255;
assign img[ 7076] = 255;
assign img[ 7077] = 255;
assign img[ 7078] = 255;
assign img[ 7079] = 255;
assign img[ 7080] = 238;
assign img[ 7081] = 254;
assign img[ 7082] = 238;
assign img[ 7083] = 255;
assign img[ 7084] = 254;
assign img[ 7085] = 255;
assign img[ 7086] = 238;
assign img[ 7087] = 223;
assign img[ 7088] = 255;
assign img[ 7089] = 255;
assign img[ 7090] = 239;
assign img[ 7091] = 206;
assign img[ 7092] = 254;
assign img[ 7093] = 255;
assign img[ 7094] = 255;
assign img[ 7095] = 255;
assign img[ 7096] = 255;
assign img[ 7097] = 255;
assign img[ 7098] = 255;
assign img[ 7099] = 255;
assign img[ 7100] = 255;
assign img[ 7101] = 255;
assign img[ 7102] = 255;
assign img[ 7103] = 255;
assign img[ 7104] = 255;
assign img[ 7105] = 255;
assign img[ 7106] = 255;
assign img[ 7107] = 255;
assign img[ 7108] = 255;
assign img[ 7109] = 255;
assign img[ 7110] = 255;
assign img[ 7111] = 255;
assign img[ 7112] = 255;
assign img[ 7113] = 255;
assign img[ 7114] = 255;
assign img[ 7115] = 255;
assign img[ 7116] = 223;
assign img[ 7117] = 239;
assign img[ 7118] = 238;
assign img[ 7119] = 238;
assign img[ 7120] = 206;
assign img[ 7121] = 238;
assign img[ 7122] = 206;
assign img[ 7123] = 236;
assign img[ 7124] = 238;
assign img[ 7125] = 238;
assign img[ 7126] = 238;
assign img[ 7127] = 238;
assign img[ 7128] = 238;
assign img[ 7129] = 254;
assign img[ 7130] = 255;
assign img[ 7131] = 255;
assign img[ 7132] = 255;
assign img[ 7133] = 255;
assign img[ 7134] = 255;
assign img[ 7135] = 223;
assign img[ 7136] = 253;
assign img[ 7137] = 255;
assign img[ 7138] = 238;
assign img[ 7139] = 238;
assign img[ 7140] = 238;
assign img[ 7141] = 255;
assign img[ 7142] = 221;
assign img[ 7143] = 238;
assign img[ 7144] = 238;
assign img[ 7145] = 255;
assign img[ 7146] = 255;
assign img[ 7147] = 239;
assign img[ 7148] = 238;
assign img[ 7149] = 238;
assign img[ 7150] = 238;
assign img[ 7151] = 223;
assign img[ 7152] = 237;
assign img[ 7153] = 255;
assign img[ 7154] = 255;
assign img[ 7155] = 255;
assign img[ 7156] = 255;
assign img[ 7157] = 255;
assign img[ 7158] = 255;
assign img[ 7159] = 255;
assign img[ 7160] = 255;
assign img[ 7161] = 191;
assign img[ 7162] = 187;
assign img[ 7163] = 187;
assign img[ 7164] = 187;
assign img[ 7165] = 255;
assign img[ 7166] = 255;
assign img[ 7167] = 255;
assign img[ 7168] = 96;
assign img[ 7169] = 206;
assign img[ 7170] = 236;
assign img[ 7171] = 238;
assign img[ 7172] = 238;
assign img[ 7173] = 254;
assign img[ 7174] = 255;
assign img[ 7175] = 255;
assign img[ 7176] = 255;
assign img[ 7177] = 255;
assign img[ 7178] = 255;
assign img[ 7179] = 255;
assign img[ 7180] = 255;
assign img[ 7181] = 255;
assign img[ 7182] = 255;
assign img[ 7183] = 223;
assign img[ 7184] = 253;
assign img[ 7185] = 238;
assign img[ 7186] = 238;
assign img[ 7187] = 206;
assign img[ 7188] = 254;
assign img[ 7189] = 255;
assign img[ 7190] = 223;
assign img[ 7191] = 255;
assign img[ 7192] = 255;
assign img[ 7193] = 255;
assign img[ 7194] = 255;
assign img[ 7195] = 255;
assign img[ 7196] = 255;
assign img[ 7197] = 255;
assign img[ 7198] = 255;
assign img[ 7199] = 207;
assign img[ 7200] = 236;
assign img[ 7201] = 254;
assign img[ 7202] = 255;
assign img[ 7203] = 255;
assign img[ 7204] = 238;
assign img[ 7205] = 255;
assign img[ 7206] = 255;
assign img[ 7207] = 255;
assign img[ 7208] = 238;
assign img[ 7209] = 238;
assign img[ 7210] = 238;
assign img[ 7211] = 238;
assign img[ 7212] = 238;
assign img[ 7213] = 238;
assign img[ 7214] = 238;
assign img[ 7215] = 238;
assign img[ 7216] = 238;
assign img[ 7217] = 238;
assign img[ 7218] = 254;
assign img[ 7219] = 255;
assign img[ 7220] = 255;
assign img[ 7221] = 255;
assign img[ 7222] = 255;
assign img[ 7223] = 255;
assign img[ 7224] = 255;
assign img[ 7225] = 255;
assign img[ 7226] = 255;
assign img[ 7227] = 255;
assign img[ 7228] = 255;
assign img[ 7229] = 255;
assign img[ 7230] = 255;
assign img[ 7231] = 255;
assign img[ 7232] = 255;
assign img[ 7233] = 255;
assign img[ 7234] = 255;
assign img[ 7235] = 255;
assign img[ 7236] = 255;
assign img[ 7237] = 191;
assign img[ 7238] = 251;
assign img[ 7239] = 255;
assign img[ 7240] = 255;
assign img[ 7241] = 255;
assign img[ 7242] = 255;
assign img[ 7243] = 239;
assign img[ 7244] = 238;
assign img[ 7245] = 238;
assign img[ 7246] = 238;
assign img[ 7247] = 238;
assign img[ 7248] = 238;
assign img[ 7249] = 255;
assign img[ 7250] = 254;
assign img[ 7251] = 255;
assign img[ 7252] = 238;
assign img[ 7253] = 238;
assign img[ 7254] = 238;
assign img[ 7255] = 238;
assign img[ 7256] = 206;
assign img[ 7257] = 254;
assign img[ 7258] = 239;
assign img[ 7259] = 239;
assign img[ 7260] = 238;
assign img[ 7261] = 255;
assign img[ 7262] = 255;
assign img[ 7263] = 255;
assign img[ 7264] = 255;
assign img[ 7265] = 239;
assign img[ 7266] = 238;
assign img[ 7267] = 238;
assign img[ 7268] = 238;
assign img[ 7269] = 238;
assign img[ 7270] = 254;
assign img[ 7271] = 255;
assign img[ 7272] = 255;
assign img[ 7273] = 239;
assign img[ 7274] = 238;
assign img[ 7275] = 238;
assign img[ 7276] = 206;
assign img[ 7277] = 238;
assign img[ 7278] = 255;
assign img[ 7279] = 239;
assign img[ 7280] = 238;
assign img[ 7281] = 238;
assign img[ 7282] = 238;
assign img[ 7283] = 238;
assign img[ 7284] = 204;
assign img[ 7285] = 236;
assign img[ 7286] = 238;
assign img[ 7287] = 238;
assign img[ 7288] = 254;
assign img[ 7289] = 255;
assign img[ 7290] = 255;
assign img[ 7291] = 255;
assign img[ 7292] = 255;
assign img[ 7293] = 255;
assign img[ 7294] = 223;
assign img[ 7295] = 255;
assign img[ 7296] = 96;
assign img[ 7297] = 239;
assign img[ 7298] = 238;
assign img[ 7299] = 238;
assign img[ 7300] = 238;
assign img[ 7301] = 239;
assign img[ 7302] = 206;
assign img[ 7303] = 204;
assign img[ 7304] = 236;
assign img[ 7305] = 238;
assign img[ 7306] = 238;
assign img[ 7307] = 254;
assign img[ 7308] = 221;
assign img[ 7309] = 221;
assign img[ 7310] = 204;
assign img[ 7311] = 206;
assign img[ 7312] = 236;
assign img[ 7313] = 238;
assign img[ 7314] = 238;
assign img[ 7315] = 238;
assign img[ 7316] = 238;
assign img[ 7317] = 238;
assign img[ 7318] = 238;
assign img[ 7319] = 238;
assign img[ 7320] = 254;
assign img[ 7321] = 255;
assign img[ 7322] = 239;
assign img[ 7323] = 255;
assign img[ 7324] = 255;
assign img[ 7325] = 255;
assign img[ 7326] = 255;
assign img[ 7327] = 255;
assign img[ 7328] = 255;
assign img[ 7329] = 255;
assign img[ 7330] = 255;
assign img[ 7331] = 255;
assign img[ 7332] = 255;
assign img[ 7333] = 207;
assign img[ 7334] = 220;
assign img[ 7335] = 221;
assign img[ 7336] = 253;
assign img[ 7337] = 223;
assign img[ 7338] = 221;
assign img[ 7339] = 253;
assign img[ 7340] = 255;
assign img[ 7341] = 239;
assign img[ 7342] = 238;
assign img[ 7343] = 238;
assign img[ 7344] = 238;
assign img[ 7345] = 239;
assign img[ 7346] = 238;
assign img[ 7347] = 238;
assign img[ 7348] = 238;
assign img[ 7349] = 238;
assign img[ 7350] = 255;
assign img[ 7351] = 255;
assign img[ 7352] = 255;
assign img[ 7353] = 255;
assign img[ 7354] = 239;
assign img[ 7355] = 254;
assign img[ 7356] = 255;
assign img[ 7357] = 223;
assign img[ 7358] = 238;
assign img[ 7359] = 255;
assign img[ 7360] = 255;
assign img[ 7361] = 255;
assign img[ 7362] = 221;
assign img[ 7363] = 253;
assign img[ 7364] = 255;
assign img[ 7365] = 255;
assign img[ 7366] = 255;
assign img[ 7367] = 255;
assign img[ 7368] = 255;
assign img[ 7369] = 239;
assign img[ 7370] = 238;
assign img[ 7371] = 238;
assign img[ 7372] = 238;
assign img[ 7373] = 238;
assign img[ 7374] = 238;
assign img[ 7375] = 238;
assign img[ 7376] = 238;
assign img[ 7377] = 238;
assign img[ 7378] = 238;
assign img[ 7379] = 254;
assign img[ 7380] = 254;
assign img[ 7381] = 223;
assign img[ 7382] = 221;
assign img[ 7383] = 253;
assign img[ 7384] = 255;
assign img[ 7385] = 255;
assign img[ 7386] = 223;
assign img[ 7387] = 255;
assign img[ 7388] = 255;
assign img[ 7389] = 255;
assign img[ 7390] = 255;
assign img[ 7391] = 255;
assign img[ 7392] = 255;
assign img[ 7393] = 239;
assign img[ 7394] = 238;
assign img[ 7395] = 238;
assign img[ 7396] = 238;
assign img[ 7397] = 255;
assign img[ 7398] = 174;
assign img[ 7399] = 170;
assign img[ 7400] = 234;
assign img[ 7401] = 255;
assign img[ 7402] = 238;
assign img[ 7403] = 239;
assign img[ 7404] = 254;
assign img[ 7405] = 254;
assign img[ 7406] = 238;
assign img[ 7407] = 222;
assign img[ 7408] = 221;
assign img[ 7409] = 221;
assign img[ 7410] = 253;
assign img[ 7411] = 239;
assign img[ 7412] = 238;
assign img[ 7413] = 255;
assign img[ 7414] = 255;
assign img[ 7415] = 255;
assign img[ 7416] = 255;
assign img[ 7417] = 255;
assign img[ 7418] = 204;
assign img[ 7419] = 238;
assign img[ 7420] = 254;
assign img[ 7421] = 255;
assign img[ 7422] = 239;
assign img[ 7423] = 238;
assign img[ 7424] = 96;
assign img[ 7425] = 206;
assign img[ 7426] = 236;
assign img[ 7427] = 238;
assign img[ 7428] = 170;
assign img[ 7429] = 170;
assign img[ 7430] = 234;
assign img[ 7431] = 238;
assign img[ 7432] = 238;
assign img[ 7433] = 254;
assign img[ 7434] = 238;
assign img[ 7435] = 238;
assign img[ 7436] = 238;
assign img[ 7437] = 238;
assign img[ 7438] = 254;
assign img[ 7439] = 255;
assign img[ 7440] = 255;
assign img[ 7441] = 255;
assign img[ 7442] = 255;
assign img[ 7443] = 191;
assign img[ 7444] = 153;
assign img[ 7445] = 253;
assign img[ 7446] = 255;
assign img[ 7447] = 255;
assign img[ 7448] = 255;
assign img[ 7449] = 255;
assign img[ 7450] = 238;
assign img[ 7451] = 238;
assign img[ 7452] = 254;
assign img[ 7453] = 255;
assign img[ 7454] = 255;
assign img[ 7455] = 223;
assign img[ 7456] = 253;
assign img[ 7457] = 255;
assign img[ 7458] = 255;
assign img[ 7459] = 255;
assign img[ 7460] = 255;
assign img[ 7461] = 255;
assign img[ 7462] = 239;
assign img[ 7463] = 238;
assign img[ 7464] = 238;
assign img[ 7465] = 238;
assign img[ 7466] = 206;
assign img[ 7467] = 206;
assign img[ 7468] = 238;
assign img[ 7469] = 255;
assign img[ 7470] = 255;
assign img[ 7471] = 255;
assign img[ 7472] = 255;
assign img[ 7473] = 255;
assign img[ 7474] = 238;
assign img[ 7475] = 238;
assign img[ 7476] = 206;
assign img[ 7477] = 254;
assign img[ 7478] = 255;
assign img[ 7479] = 255;
assign img[ 7480] = 238;
assign img[ 7481] = 255;
assign img[ 7482] = 255;
assign img[ 7483] = 255;
assign img[ 7484] = 255;
assign img[ 7485] = 255;
assign img[ 7486] = 255;
assign img[ 7487] = 255;
assign img[ 7488] = 255;
assign img[ 7489] = 255;
assign img[ 7490] = 255;
assign img[ 7491] = 255;
assign img[ 7492] = 255;
assign img[ 7493] = 239;
assign img[ 7494] = 238;
assign img[ 7495] = 238;
assign img[ 7496] = 238;
assign img[ 7497] = 238;
assign img[ 7498] = 254;
assign img[ 7499] = 223;
assign img[ 7500] = 221;
assign img[ 7501] = 255;
assign img[ 7502] = 238;
assign img[ 7503] = 254;
assign img[ 7504] = 255;
assign img[ 7505] = 255;
assign img[ 7506] = 238;
assign img[ 7507] = 255;
assign img[ 7508] = 223;
assign img[ 7509] = 223;
assign img[ 7510] = 255;
assign img[ 7511] = 255;
assign img[ 7512] = 239;
assign img[ 7513] = 238;
assign img[ 7514] = 238;
assign img[ 7515] = 238;
assign img[ 7516] = 254;
assign img[ 7517] = 255;
assign img[ 7518] = 255;
assign img[ 7519] = 239;
assign img[ 7520] = 238;
assign img[ 7521] = 238;
assign img[ 7522] = 238;
assign img[ 7523] = 238;
assign img[ 7524] = 238;
assign img[ 7525] = 239;
assign img[ 7526] = 238;
assign img[ 7527] = 238;
assign img[ 7528] = 238;
assign img[ 7529] = 255;
assign img[ 7530] = 255;
assign img[ 7531] = 239;
assign img[ 7532] = 238;
assign img[ 7533] = 255;
assign img[ 7534] = 223;
assign img[ 7535] = 253;
assign img[ 7536] = 255;
assign img[ 7537] = 255;
assign img[ 7538] = 255;
assign img[ 7539] = 239;
assign img[ 7540] = 254;
assign img[ 7541] = 255;
assign img[ 7542] = 254;
assign img[ 7543] = 255;
assign img[ 7544] = 254;
assign img[ 7545] = 255;
assign img[ 7546] = 255;
assign img[ 7547] = 255;
assign img[ 7548] = 255;
assign img[ 7549] = 255;
assign img[ 7550] = 223;
assign img[ 7551] = 255;
assign img[ 7552] = 96;
assign img[ 7553] = 206;
assign img[ 7554] = 252;
assign img[ 7555] = 255;
assign img[ 7556] = 223;
assign img[ 7557] = 253;
assign img[ 7558] = 191;
assign img[ 7559] = 187;
assign img[ 7560] = 251;
assign img[ 7561] = 255;
assign img[ 7562] = 254;
assign img[ 7563] = 223;
assign img[ 7564] = 205;
assign img[ 7565] = 204;
assign img[ 7566] = 236;
assign img[ 7567] = 207;
assign img[ 7568] = 252;
assign img[ 7569] = 238;
assign img[ 7570] = 238;
assign img[ 7571] = 239;
assign img[ 7572] = 254;
assign img[ 7573] = 255;
assign img[ 7574] = 239;
assign img[ 7575] = 238;
assign img[ 7576] = 238;
assign img[ 7577] = 238;
assign img[ 7578] = 238;
assign img[ 7579] = 238;
assign img[ 7580] = 238;
assign img[ 7581] = 238;
assign img[ 7582] = 238;
assign img[ 7583] = 142;
assign img[ 7584] = 236;
assign img[ 7585] = 238;
assign img[ 7586] = 238;
assign img[ 7587] = 238;
assign img[ 7588] = 255;
assign img[ 7589] = 255;
assign img[ 7590] = 255;
assign img[ 7591] = 255;
assign img[ 7592] = 255;
assign img[ 7593] = 255;
assign img[ 7594] = 255;
assign img[ 7595] = 255;
assign img[ 7596] = 255;
assign img[ 7597] = 255;
assign img[ 7598] = 255;
assign img[ 7599] = 255;
assign img[ 7600] = 254;
assign img[ 7601] = 255;
assign img[ 7602] = 254;
assign img[ 7603] = 255;
assign img[ 7604] = 221;
assign img[ 7605] = 253;
assign img[ 7606] = 255;
assign img[ 7607] = 255;
assign img[ 7608] = 239;
assign img[ 7609] = 255;
assign img[ 7610] = 255;
assign img[ 7611] = 255;
assign img[ 7612] = 255;
assign img[ 7613] = 255;
assign img[ 7614] = 255;
assign img[ 7615] = 255;
assign img[ 7616] = 255;
assign img[ 7617] = 255;
assign img[ 7618] = 255;
assign img[ 7619] = 255;
assign img[ 7620] = 255;
assign img[ 7621] = 239;
assign img[ 7622] = 254;
assign img[ 7623] = 239;
assign img[ 7624] = 238;
assign img[ 7625] = 238;
assign img[ 7626] = 254;
assign img[ 7627] = 223;
assign img[ 7628] = 255;
assign img[ 7629] = 255;
assign img[ 7630] = 254;
assign img[ 7631] = 255;
assign img[ 7632] = 254;
assign img[ 7633] = 255;
assign img[ 7634] = 255;
assign img[ 7635] = 255;
assign img[ 7636] = 255;
assign img[ 7637] = 239;
assign img[ 7638] = 238;
assign img[ 7639] = 238;
assign img[ 7640] = 238;
assign img[ 7641] = 238;
assign img[ 7642] = 238;
assign img[ 7643] = 238;
assign img[ 7644] = 238;
assign img[ 7645] = 255;
assign img[ 7646] = 254;
assign img[ 7647] = 255;
assign img[ 7648] = 155;
assign img[ 7649] = 217;
assign img[ 7650] = 236;
assign img[ 7651] = 238;
assign img[ 7652] = 238;
assign img[ 7653] = 238;
assign img[ 7654] = 238;
assign img[ 7655] = 238;
assign img[ 7656] = 238;
assign img[ 7657] = 255;
assign img[ 7658] = 255;
assign img[ 7659] = 175;
assign img[ 7660] = 170;
assign img[ 7661] = 238;
assign img[ 7662] = 238;
assign img[ 7663] = 238;
assign img[ 7664] = 238;
assign img[ 7665] = 238;
assign img[ 7666] = 238;
assign img[ 7667] = 238;
assign img[ 7668] = 206;
assign img[ 7669] = 255;
assign img[ 7670] = 255;
assign img[ 7671] = 255;
assign img[ 7672] = 255;
assign img[ 7673] = 255;
assign img[ 7674] = 238;
assign img[ 7675] = 238;
assign img[ 7676] = 220;
assign img[ 7677] = 255;
assign img[ 7678] = 255;
assign img[ 7679] = 255;
assign img[ 7680] = 64;
assign img[ 7681] = 68;
assign img[ 7682] = 116;
assign img[ 7683] = 255;
assign img[ 7684] = 255;
assign img[ 7685] = 255;
assign img[ 7686] = 238;
assign img[ 7687] = 238;
assign img[ 7688] = 238;
assign img[ 7689] = 238;
assign img[ 7690] = 238;
assign img[ 7691] = 238;
assign img[ 7692] = 187;
assign img[ 7693] = 251;
assign img[ 7694] = 255;
assign img[ 7695] = 255;
assign img[ 7696] = 205;
assign img[ 7697] = 204;
assign img[ 7698] = 236;
assign img[ 7699] = 238;
assign img[ 7700] = 238;
assign img[ 7701] = 238;
assign img[ 7702] = 238;
assign img[ 7703] = 238;
assign img[ 7704] = 238;
assign img[ 7705] = 255;
assign img[ 7706] = 255;
assign img[ 7707] = 255;
assign img[ 7708] = 238;
assign img[ 7709] = 238;
assign img[ 7710] = 238;
assign img[ 7711] = 238;
assign img[ 7712] = 238;
assign img[ 7713] = 238;
assign img[ 7714] = 238;
assign img[ 7715] = 255;
assign img[ 7716] = 255;
assign img[ 7717] = 255;
assign img[ 7718] = 255;
assign img[ 7719] = 255;
assign img[ 7720] = 255;
assign img[ 7721] = 255;
assign img[ 7722] = 255;
assign img[ 7723] = 255;
assign img[ 7724] = 255;
assign img[ 7725] = 255;
assign img[ 7726] = 238;
assign img[ 7727] = 255;
assign img[ 7728] = 255;
assign img[ 7729] = 255;
assign img[ 7730] = 255;
assign img[ 7731] = 255;
assign img[ 7732] = 255;
assign img[ 7733] = 255;
assign img[ 7734] = 255;
assign img[ 7735] = 255;
assign img[ 7736] = 255;
assign img[ 7737] = 255;
assign img[ 7738] = 239;
assign img[ 7739] = 238;
assign img[ 7740] = 238;
assign img[ 7741] = 223;
assign img[ 7742] = 221;
assign img[ 7743] = 255;
assign img[ 7744] = 255;
assign img[ 7745] = 255;
assign img[ 7746] = 255;
assign img[ 7747] = 255;
assign img[ 7748] = 255;
assign img[ 7749] = 239;
assign img[ 7750] = 238;
assign img[ 7751] = 238;
assign img[ 7752] = 238;
assign img[ 7753] = 238;
assign img[ 7754] = 238;
assign img[ 7755] = 254;
assign img[ 7756] = 254;
assign img[ 7757] = 255;
assign img[ 7758] = 255;
assign img[ 7759] = 255;
assign img[ 7760] = 223;
assign img[ 7761] = 255;
assign img[ 7762] = 223;
assign img[ 7763] = 253;
assign img[ 7764] = 255;
assign img[ 7765] = 255;
assign img[ 7766] = 238;
assign img[ 7767] = 255;
assign img[ 7768] = 222;
assign img[ 7769] = 255;
assign img[ 7770] = 255;
assign img[ 7771] = 255;
assign img[ 7772] = 255;
assign img[ 7773] = 255;
assign img[ 7774] = 255;
assign img[ 7775] = 255;
assign img[ 7776] = 191;
assign img[ 7777] = 187;
assign img[ 7778] = 234;
assign img[ 7779] = 254;
assign img[ 7780] = 238;
assign img[ 7781] = 238;
assign img[ 7782] = 204;
assign img[ 7783] = 238;
assign img[ 7784] = 238;
assign img[ 7785] = 238;
assign img[ 7786] = 238;
assign img[ 7787] = 255;
assign img[ 7788] = 255;
assign img[ 7789] = 255;
assign img[ 7790] = 223;
assign img[ 7791] = 221;
assign img[ 7792] = 204;
assign img[ 7793] = 252;
assign img[ 7794] = 255;
assign img[ 7795] = 255;
assign img[ 7796] = 221;
assign img[ 7797] = 255;
assign img[ 7798] = 255;
assign img[ 7799] = 255;
assign img[ 7800] = 255;
assign img[ 7801] = 239;
assign img[ 7802] = 238;
assign img[ 7803] = 255;
assign img[ 7804] = 255;
assign img[ 7805] = 255;
assign img[ 7806] = 207;
assign img[ 7807] = 204;
assign img[ 7808] = 64;
assign img[ 7809] = 68;
assign img[ 7810] = 100;
assign img[ 7811] = 238;
assign img[ 7812] = 254;
assign img[ 7813] = 239;
assign img[ 7814] = 238;
assign img[ 7815] = 238;
assign img[ 7816] = 238;
assign img[ 7817] = 255;
assign img[ 7818] = 204;
assign img[ 7819] = 238;
assign img[ 7820] = 238;
assign img[ 7821] = 221;
assign img[ 7822] = 221;
assign img[ 7823] = 205;
assign img[ 7824] = 204;
assign img[ 7825] = 236;
assign img[ 7826] = 238;
assign img[ 7827] = 174;
assign img[ 7828] = 170;
assign img[ 7829] = 238;
assign img[ 7830] = 254;
assign img[ 7831] = 255;
assign img[ 7832] = 255;
assign img[ 7833] = 255;
assign img[ 7834] = 187;
assign img[ 7835] = 255;
assign img[ 7836] = 255;
assign img[ 7837] = 255;
assign img[ 7838] = 255;
assign img[ 7839] = 255;
assign img[ 7840] = 238;
assign img[ 7841] = 238;
assign img[ 7842] = 238;
assign img[ 7843] = 238;
assign img[ 7844] = 238;
assign img[ 7845] = 238;
assign img[ 7846] = 204;
assign img[ 7847] = 238;
assign img[ 7848] = 238;
assign img[ 7849] = 238;
assign img[ 7850] = 254;
assign img[ 7851] = 255;
assign img[ 7852] = 255;
assign img[ 7853] = 255;
assign img[ 7854] = 255;
assign img[ 7855] = 255;
assign img[ 7856] = 255;
assign img[ 7857] = 255;
assign img[ 7858] = 255;
assign img[ 7859] = 239;
assign img[ 7860] = 238;
assign img[ 7861] = 254;
assign img[ 7862] = 239;
assign img[ 7863] = 255;
assign img[ 7864] = 255;
assign img[ 7865] = 239;
assign img[ 7866] = 204;
assign img[ 7867] = 238;
assign img[ 7868] = 238;
assign img[ 7869] = 223;
assign img[ 7870] = 236;
assign img[ 7871] = 238;
assign img[ 7872] = 238;
assign img[ 7873] = 191;
assign img[ 7874] = 139;
assign img[ 7875] = 238;
assign img[ 7876] = 238;
assign img[ 7877] = 238;
assign img[ 7878] = 238;
assign img[ 7879] = 238;
assign img[ 7880] = 238;
assign img[ 7881] = 238;
assign img[ 7882] = 254;
assign img[ 7883] = 255;
assign img[ 7884] = 221;
assign img[ 7885] = 255;
assign img[ 7886] = 255;
assign img[ 7887] = 255;
assign img[ 7888] = 255;
assign img[ 7889] = 255;
assign img[ 7890] = 255;
assign img[ 7891] = 255;
assign img[ 7892] = 255;
assign img[ 7893] = 255;
assign img[ 7894] = 238;
assign img[ 7895] = 238;
assign img[ 7896] = 223;
assign img[ 7897] = 221;
assign img[ 7898] = 221;
assign img[ 7899] = 237;
assign img[ 7900] = 238;
assign img[ 7901] = 238;
assign img[ 7902] = 254;
assign img[ 7903] = 255;
assign img[ 7904] = 238;
assign img[ 7905] = 238;
assign img[ 7906] = 254;
assign img[ 7907] = 255;
assign img[ 7908] = 255;
assign img[ 7909] = 255;
assign img[ 7910] = 157;
assign img[ 7911] = 255;
assign img[ 7912] = 255;
assign img[ 7913] = 255;
assign img[ 7914] = 238;
assign img[ 7915] = 238;
assign img[ 7916] = 254;
assign img[ 7917] = 255;
assign img[ 7918] = 255;
assign img[ 7919] = 255;
assign img[ 7920] = 255;
assign img[ 7921] = 223;
assign img[ 7922] = 221;
assign img[ 7923] = 223;
assign img[ 7924] = 255;
assign img[ 7925] = 255;
assign img[ 7926] = 207;
assign img[ 7927] = 236;
assign img[ 7928] = 254;
assign img[ 7929] = 207;
assign img[ 7930] = 204;
assign img[ 7931] = 206;
assign img[ 7932] = 221;
assign img[ 7933] = 221;
assign img[ 7934] = 221;
assign img[ 7935] = 221;
assign img[ 7936] = 96;
assign img[ 7937] = 206;
assign img[ 7938] = 236;
assign img[ 7939] = 238;
assign img[ 7940] = 255;
assign img[ 7941] = 255;
assign img[ 7942] = 223;
assign img[ 7943] = 221;
assign img[ 7944] = 253;
assign img[ 7945] = 255;
assign img[ 7946] = 255;
assign img[ 7947] = 255;
assign img[ 7948] = 239;
assign img[ 7949] = 238;
assign img[ 7950] = 238;
assign img[ 7951] = 238;
assign img[ 7952] = 238;
assign img[ 7953] = 238;
assign img[ 7954] = 238;
assign img[ 7955] = 238;
assign img[ 7956] = 238;
assign img[ 7957] = 254;
assign img[ 7958] = 155;
assign img[ 7959] = 255;
assign img[ 7960] = 255;
assign img[ 7961] = 255;
assign img[ 7962] = 207;
assign img[ 7963] = 238;
assign img[ 7964] = 238;
assign img[ 7965] = 238;
assign img[ 7966] = 238;
assign img[ 7967] = 255;
assign img[ 7968] = 255;
assign img[ 7969] = 255;
assign img[ 7970] = 238;
assign img[ 7971] = 255;
assign img[ 7972] = 239;
assign img[ 7973] = 238;
assign img[ 7974] = 254;
assign img[ 7975] = 255;
assign img[ 7976] = 255;
assign img[ 7977] = 255;
assign img[ 7978] = 238;
assign img[ 7979] = 238;
assign img[ 7980] = 238;
assign img[ 7981] = 238;
assign img[ 7982] = 238;
assign img[ 7983] = 255;
assign img[ 7984] = 255;
assign img[ 7985] = 255;
assign img[ 7986] = 255;
assign img[ 7987] = 255;
assign img[ 7988] = 255;
assign img[ 7989] = 255;
assign img[ 7990] = 255;
assign img[ 7991] = 255;
assign img[ 7992] = 255;
assign img[ 7993] = 255;
assign img[ 7994] = 255;
assign img[ 7995] = 239;
assign img[ 7996] = 238;
assign img[ 7997] = 238;
assign img[ 7998] = 254;
assign img[ 7999] = 255;
assign img[ 8000] = 255;
assign img[ 8001] = 255;
assign img[ 8002] = 255;
assign img[ 8003] = 255;
assign img[ 8004] = 255;
assign img[ 8005] = 255;
assign img[ 8006] = 255;
assign img[ 8007] = 255;
assign img[ 8008] = 255;
assign img[ 8009] = 255;
assign img[ 8010] = 255;
assign img[ 8011] = 255;
assign img[ 8012] = 238;
assign img[ 8013] = 238;
assign img[ 8014] = 238;
assign img[ 8015] = 255;
assign img[ 8016] = 255;
assign img[ 8017] = 255;
assign img[ 8018] = 255;
assign img[ 8019] = 255;
assign img[ 8020] = 255;
assign img[ 8021] = 255;
assign img[ 8022] = 238;
assign img[ 8023] = 238;
assign img[ 8024] = 254;
assign img[ 8025] = 255;
assign img[ 8026] = 255;
assign img[ 8027] = 255;
assign img[ 8028] = 255;
assign img[ 8029] = 255;
assign img[ 8030] = 239;
assign img[ 8031] = 238;
assign img[ 8032] = 238;
assign img[ 8033] = 238;
assign img[ 8034] = 238;
assign img[ 8035] = 238;
assign img[ 8036] = 238;
assign img[ 8037] = 255;
assign img[ 8038] = 204;
assign img[ 8039] = 238;
assign img[ 8040] = 254;
assign img[ 8041] = 239;
assign img[ 8042] = 238;
assign img[ 8043] = 238;
assign img[ 8044] = 254;
assign img[ 8045] = 239;
assign img[ 8046] = 238;
assign img[ 8047] = 238;
assign img[ 8048] = 238;
assign img[ 8049] = 254;
assign img[ 8050] = 238;
assign img[ 8051] = 238;
assign img[ 8052] = 238;
assign img[ 8053] = 238;
assign img[ 8054] = 238;
assign img[ 8055] = 254;
assign img[ 8056] = 238;
assign img[ 8057] = 238;
assign img[ 8058] = 220;
assign img[ 8059] = 255;
assign img[ 8060] = 255;
assign img[ 8061] = 255;
assign img[ 8062] = 223;
assign img[ 8063] = 255;
assign img[ 8064] = 64;
assign img[ 8065] = 132;
assign img[ 8066] = 216;
assign img[ 8067] = 205;
assign img[ 8068] = 204;
assign img[ 8069] = 204;
assign img[ 8070] = 190;
assign img[ 8071] = 255;
assign img[ 8072] = 255;
assign img[ 8073] = 255;
assign img[ 8074] = 255;
assign img[ 8075] = 255;
assign img[ 8076] = 191;
assign img[ 8077] = 155;
assign img[ 8078] = 153;
assign img[ 8079] = 153;
assign img[ 8080] = 217;
assign img[ 8081] = 221;
assign img[ 8082] = 253;
assign img[ 8083] = 255;
assign img[ 8084] = 255;
assign img[ 8085] = 255;
assign img[ 8086] = 255;
assign img[ 8087] = 255;
assign img[ 8088] = 255;
assign img[ 8089] = 255;
assign img[ 8090] = 239;
assign img[ 8091] = 238;
assign img[ 8092] = 238;
assign img[ 8093] = 255;
assign img[ 8094] = 255;
assign img[ 8095] = 255;
assign img[ 8096] = 255;
assign img[ 8097] = 255;
assign img[ 8098] = 255;
assign img[ 8099] = 255;
assign img[ 8100] = 255;
assign img[ 8101] = 255;
assign img[ 8102] = 238;
assign img[ 8103] = 238;
assign img[ 8104] = 238;
assign img[ 8105] = 255;
assign img[ 8106] = 255;
assign img[ 8107] = 255;
assign img[ 8108] = 254;
assign img[ 8109] = 255;
assign img[ 8110] = 255;
assign img[ 8111] = 223;
assign img[ 8112] = 255;
assign img[ 8113] = 255;
assign img[ 8114] = 255;
assign img[ 8115] = 255;
assign img[ 8116] = 255;
assign img[ 8117] = 255;
assign img[ 8118] = 255;
assign img[ 8119] = 255;
assign img[ 8120] = 255;
assign img[ 8121] = 255;
assign img[ 8122] = 255;
assign img[ 8123] = 255;
assign img[ 8124] = 255;
assign img[ 8125] = 255;
assign img[ 8126] = 238;
assign img[ 8127] = 255;
assign img[ 8128] = 255;
assign img[ 8129] = 255;
assign img[ 8130] = 239;
assign img[ 8131] = 238;
assign img[ 8132] = 238;
assign img[ 8133] = 238;
assign img[ 8134] = 254;
assign img[ 8135] = 255;
assign img[ 8136] = 255;
assign img[ 8137] = 255;
assign img[ 8138] = 255;
assign img[ 8139] = 255;
assign img[ 8140] = 255;
assign img[ 8141] = 255;
assign img[ 8142] = 255;
assign img[ 8143] = 255;
assign img[ 8144] = 223;
assign img[ 8145] = 255;
assign img[ 8146] = 255;
assign img[ 8147] = 255;
assign img[ 8148] = 255;
assign img[ 8149] = 239;
assign img[ 8150] = 238;
assign img[ 8151] = 238;
assign img[ 8152] = 222;
assign img[ 8153] = 255;
assign img[ 8154] = 239;
assign img[ 8155] = 238;
assign img[ 8156] = 254;
assign img[ 8157] = 255;
assign img[ 8158] = 255;
assign img[ 8159] = 255;
assign img[ 8160] = 255;
assign img[ 8161] = 239;
assign img[ 8162] = 254;
assign img[ 8163] = 255;
assign img[ 8164] = 255;
assign img[ 8165] = 239;
assign img[ 8166] = 174;
assign img[ 8167] = 239;
assign img[ 8168] = 255;
assign img[ 8169] = 239;
assign img[ 8170] = 238;
assign img[ 8171] = 238;
assign img[ 8172] = 204;
assign img[ 8173] = 255;
assign img[ 8174] = 255;
assign img[ 8175] = 255;
assign img[ 8176] = 255;
assign img[ 8177] = 255;
assign img[ 8178] = 223;
assign img[ 8179] = 191;
assign img[ 8180] = 187;
assign img[ 8181] = 255;
assign img[ 8182] = 255;
assign img[ 8183] = 255;
assign img[ 8184] = 255;
assign img[ 8185] = 255;
assign img[ 8186] = 171;
assign img[ 8187] = 234;
assign img[ 8188] = 234;
assign img[ 8189] = 234;
assign img[ 8190] = 186;
assign img[ 8191] = 235;
assign img[ 8192] = 16;
assign img[ 8193] = 221;
assign img[ 8194] = 253;
assign img[ 8195] = 223;
assign img[ 8196] = 205;
assign img[ 8197] = 204;
assign img[ 8198] = 236;
assign img[ 8199] = 238;
assign img[ 8200] = 238;
assign img[ 8201] = 238;
assign img[ 8202] = 238;
assign img[ 8203] = 238;
assign img[ 8204] = 238;
assign img[ 8205] = 238;
assign img[ 8206] = 204;
assign img[ 8207] = 238;
assign img[ 8208] = 238;
assign img[ 8209] = 255;
assign img[ 8210] = 255;
assign img[ 8211] = 223;
assign img[ 8212] = 236;
assign img[ 8213] = 239;
assign img[ 8214] = 255;
assign img[ 8215] = 223;
assign img[ 8216] = 236;
assign img[ 8217] = 191;
assign img[ 8218] = 187;
assign img[ 8219] = 255;
assign img[ 8220] = 255;
assign img[ 8221] = 255;
assign img[ 8222] = 255;
assign img[ 8223] = 191;
assign img[ 8224] = 170;
assign img[ 8225] = 251;
assign img[ 8226] = 255;
assign img[ 8227] = 255;
assign img[ 8228] = 255;
assign img[ 8229] = 239;
assign img[ 8230] = 238;
assign img[ 8231] = 238;
assign img[ 8232] = 238;
assign img[ 8233] = 238;
assign img[ 8234] = 254;
assign img[ 8235] = 255;
assign img[ 8236] = 239;
assign img[ 8237] = 254;
assign img[ 8238] = 207;
assign img[ 8239] = 204;
assign img[ 8240] = 236;
assign img[ 8241] = 238;
assign img[ 8242] = 238;
assign img[ 8243] = 255;
assign img[ 8244] = 238;
assign img[ 8245] = 238;
assign img[ 8246] = 206;
assign img[ 8247] = 206;
assign img[ 8248] = 238;
assign img[ 8249] = 238;
assign img[ 8250] = 222;
assign img[ 8251] = 255;
assign img[ 8252] = 255;
assign img[ 8253] = 159;
assign img[ 8254] = 255;
assign img[ 8255] = 255;
assign img[ 8256] = 255;
assign img[ 8257] = 255;
assign img[ 8258] = 191;
assign img[ 8259] = 255;
assign img[ 8260] = 255;
assign img[ 8261] = 255;
assign img[ 8262] = 255;
assign img[ 8263] = 255;
assign img[ 8264] = 239;
assign img[ 8265] = 206;
assign img[ 8266] = 236;
assign img[ 8267] = 239;
assign img[ 8268] = 238;
assign img[ 8269] = 254;
assign img[ 8270] = 255;
assign img[ 8271] = 239;
assign img[ 8272] = 255;
assign img[ 8273] = 255;
assign img[ 8274] = 238;
assign img[ 8275] = 238;
assign img[ 8276] = 238;
assign img[ 8277] = 238;
assign img[ 8278] = 238;
assign img[ 8279] = 238;
assign img[ 8280] = 254;
assign img[ 8281] = 255;
assign img[ 8282] = 255;
assign img[ 8283] = 255;
assign img[ 8284] = 255;
assign img[ 8285] = 255;
assign img[ 8286] = 255;
assign img[ 8287] = 191;
assign img[ 8288] = 171;
assign img[ 8289] = 170;
assign img[ 8290] = 250;
assign img[ 8291] = 255;
assign img[ 8292] = 255;
assign img[ 8293] = 255;
assign img[ 8294] = 238;
assign img[ 8295] = 255;
assign img[ 8296] = 238;
assign img[ 8297] = 206;
assign img[ 8298] = 236;
assign img[ 8299] = 238;
assign img[ 8300] = 222;
assign img[ 8301] = 255;
assign img[ 8302] = 223;
assign img[ 8303] = 205;
assign img[ 8304] = 220;
assign img[ 8305] = 221;
assign img[ 8306] = 221;
assign img[ 8307] = 221;
assign img[ 8308] = 221;
assign img[ 8309] = 205;
assign img[ 8310] = 238;
assign img[ 8311] = 238;
assign img[ 8312] = 238;
assign img[ 8313] = 255;
assign img[ 8314] = 255;
assign img[ 8315] = 223;
assign img[ 8316] = 221;
assign img[ 8317] = 253;
assign img[ 8318] = 207;
assign img[ 8319] = 238;
assign img[ 8320] = 80;
assign img[ 8321] = 85;
assign img[ 8322] = 117;
assign img[ 8323] = 206;
assign img[ 8324] = 204;
assign img[ 8325] = 204;
assign img[ 8326] = 220;
assign img[ 8327] = 221;
assign img[ 8328] = 253;
assign img[ 8329] = 239;
assign img[ 8330] = 254;
assign img[ 8331] = 255;
assign img[ 8332] = 255;
assign img[ 8333] = 255;
assign img[ 8334] = 255;
assign img[ 8335] = 239;
assign img[ 8336] = 254;
assign img[ 8337] = 239;
assign img[ 8338] = 254;
assign img[ 8339] = 239;
assign img[ 8340] = 204;
assign img[ 8341] = 238;
assign img[ 8342] = 206;
assign img[ 8343] = 254;
assign img[ 8344] = 255;
assign img[ 8345] = 191;
assign img[ 8346] = 251;
assign img[ 8347] = 255;
assign img[ 8348] = 255;
assign img[ 8349] = 255;
assign img[ 8350] = 255;
assign img[ 8351] = 191;
assign img[ 8352] = 187;
assign img[ 8353] = 251;
assign img[ 8354] = 255;
assign img[ 8355] = 255;
assign img[ 8356] = 239;
assign img[ 8357] = 255;
assign img[ 8358] = 255;
assign img[ 8359] = 255;
assign img[ 8360] = 255;
assign img[ 8361] = 255;
assign img[ 8362] = 255;
assign img[ 8363] = 255;
assign img[ 8364] = 207;
assign img[ 8365] = 204;
assign img[ 8366] = 236;
assign img[ 8367] = 255;
assign img[ 8368] = 255;
assign img[ 8369] = 255;
assign img[ 8370] = 255;
assign img[ 8371] = 223;
assign img[ 8372] = 221;
assign img[ 8373] = 255;
assign img[ 8374] = 255;
assign img[ 8375] = 255;
assign img[ 8376] = 255;
assign img[ 8377] = 255;
assign img[ 8378] = 223;
assign img[ 8379] = 255;
assign img[ 8380] = 255;
assign img[ 8381] = 255;
assign img[ 8382] = 238;
assign img[ 8383] = 238;
assign img[ 8384] = 238;
assign img[ 8385] = 255;
assign img[ 8386] = 238;
assign img[ 8387] = 238;
assign img[ 8388] = 238;
assign img[ 8389] = 238;
assign img[ 8390] = 254;
assign img[ 8391] = 255;
assign img[ 8392] = 238;
assign img[ 8393] = 238;
assign img[ 8394] = 254;
assign img[ 8395] = 239;
assign img[ 8396] = 238;
assign img[ 8397] = 238;
assign img[ 8398] = 238;
assign img[ 8399] = 255;
assign img[ 8400] = 239;
assign img[ 8401] = 238;
assign img[ 8402] = 206;
assign img[ 8403] = 207;
assign img[ 8404] = 204;
assign img[ 8405] = 239;
assign img[ 8406] = 238;
assign img[ 8407] = 238;
assign img[ 8408] = 238;
assign img[ 8409] = 238;
assign img[ 8410] = 238;
assign img[ 8411] = 255;
assign img[ 8412] = 255;
assign img[ 8413] = 239;
assign img[ 8414] = 254;
assign img[ 8415] = 255;
assign img[ 8416] = 170;
assign img[ 8417] = 234;
assign img[ 8418] = 255;
assign img[ 8419] = 255;
assign img[ 8420] = 238;
assign img[ 8421] = 238;
assign img[ 8422] = 238;
assign img[ 8423] = 238;
assign img[ 8424] = 255;
assign img[ 8425] = 255;
assign img[ 8426] = 238;
assign img[ 8427] = 255;
assign img[ 8428] = 238;
assign img[ 8429] = 238;
assign img[ 8430] = 204;
assign img[ 8431] = 204;
assign img[ 8432] = 204;
assign img[ 8433] = 221;
assign img[ 8434] = 255;
assign img[ 8435] = 255;
assign img[ 8436] = 238;
assign img[ 8437] = 238;
assign img[ 8438] = 238;
assign img[ 8439] = 238;
assign img[ 8440] = 238;
assign img[ 8441] = 238;
assign img[ 8442] = 170;
assign img[ 8443] = 170;
assign img[ 8444] = 206;
assign img[ 8445] = 238;
assign img[ 8446] = 206;
assign img[ 8447] = 204;
assign img[ 8448] = 96;
assign img[ 8449] = 223;
assign img[ 8450] = 205;
assign img[ 8451] = 204;
assign img[ 8452] = 172;
assign img[ 8453] = 186;
assign img[ 8454] = 139;
assign img[ 8455] = 238;
assign img[ 8456] = 238;
assign img[ 8457] = 239;
assign img[ 8458] = 238;
assign img[ 8459] = 255;
assign img[ 8460] = 239;
assign img[ 8461] = 238;
assign img[ 8462] = 254;
assign img[ 8463] = 223;
assign img[ 8464] = 204;
assign img[ 8465] = 204;
assign img[ 8466] = 236;
assign img[ 8467] = 239;
assign img[ 8468] = 238;
assign img[ 8469] = 238;
assign img[ 8470] = 238;
assign img[ 8471] = 239;
assign img[ 8472] = 238;
assign img[ 8473] = 238;
assign img[ 8474] = 220;
assign img[ 8475] = 255;
assign img[ 8476] = 255;
assign img[ 8477] = 255;
assign img[ 8478] = 255;
assign img[ 8479] = 191;
assign img[ 8480] = 255;
assign img[ 8481] = 255;
assign img[ 8482] = 238;
assign img[ 8483] = 255;
assign img[ 8484] = 254;
assign img[ 8485] = 255;
assign img[ 8486] = 255;
assign img[ 8487] = 191;
assign img[ 8488] = 255;
assign img[ 8489] = 255;
assign img[ 8490] = 255;
assign img[ 8491] = 255;
assign img[ 8492] = 255;
assign img[ 8493] = 255;
assign img[ 8494] = 255;
assign img[ 8495] = 223;
assign img[ 8496] = 255;
assign img[ 8497] = 255;
assign img[ 8498] = 255;
assign img[ 8499] = 255;
assign img[ 8500] = 255;
assign img[ 8501] = 255;
assign img[ 8502] = 255;
assign img[ 8503] = 255;
assign img[ 8504] = 255;
assign img[ 8505] = 255;
assign img[ 8506] = 255;
assign img[ 8507] = 255;
assign img[ 8508] = 255;
assign img[ 8509] = 255;
assign img[ 8510] = 223;
assign img[ 8511] = 255;
assign img[ 8512] = 255;
assign img[ 8513] = 239;
assign img[ 8514] = 204;
assign img[ 8515] = 238;
assign img[ 8516] = 254;
assign img[ 8517] = 223;
assign img[ 8518] = 255;
assign img[ 8519] = 255;
assign img[ 8520] = 254;
assign img[ 8521] = 255;
assign img[ 8522] = 255;
assign img[ 8523] = 239;
assign img[ 8524] = 238;
assign img[ 8525] = 238;
assign img[ 8526] = 238;
assign img[ 8527] = 255;
assign img[ 8528] = 255;
assign img[ 8529] = 255;
assign img[ 8530] = 223;
assign img[ 8531] = 255;
assign img[ 8532] = 255;
assign img[ 8533] = 239;
assign img[ 8534] = 238;
assign img[ 8535] = 238;
assign img[ 8536] = 190;
assign img[ 8537] = 187;
assign img[ 8538] = 251;
assign img[ 8539] = 255;
assign img[ 8540] = 255;
assign img[ 8541] = 255;
assign img[ 8542] = 255;
assign img[ 8543] = 191;
assign img[ 8544] = 187;
assign img[ 8545] = 251;
assign img[ 8546] = 255;
assign img[ 8547] = 255;
assign img[ 8548] = 255;
assign img[ 8549] = 255;
assign img[ 8550] = 187;
assign img[ 8551] = 187;
assign img[ 8552] = 255;
assign img[ 8553] = 255;
assign img[ 8554] = 255;
assign img[ 8555] = 255;
assign img[ 8556] = 239;
assign img[ 8557] = 238;
assign img[ 8558] = 238;
assign img[ 8559] = 238;
assign img[ 8560] = 238;
assign img[ 8561] = 238;
assign img[ 8562] = 238;
assign img[ 8563] = 255;
assign img[ 8564] = 255;
assign img[ 8565] = 255;
assign img[ 8566] = 239;
assign img[ 8567] = 238;
assign img[ 8568] = 238;
assign img[ 8569] = 207;
assign img[ 8570] = 204;
assign img[ 8571] = 141;
assign img[ 8572] = 236;
assign img[ 8573] = 238;
assign img[ 8574] = 238;
assign img[ 8575] = 238;
assign img[ 8576] = 96;
assign img[ 8577] = 238;
assign img[ 8578] = 238;
assign img[ 8579] = 207;
assign img[ 8580] = 204;
assign img[ 8581] = 236;
assign img[ 8582] = 174;
assign img[ 8583] = 186;
assign img[ 8584] = 251;
assign img[ 8585] = 255;
assign img[ 8586] = 238;
assign img[ 8587] = 238;
assign img[ 8588] = 238;
assign img[ 8589] = 238;
assign img[ 8590] = 238;
assign img[ 8591] = 238;
assign img[ 8592] = 204;
assign img[ 8593] = 236;
assign img[ 8594] = 255;
assign img[ 8595] = 255;
assign img[ 8596] = 238;
assign img[ 8597] = 238;
assign img[ 8598] = 238;
assign img[ 8599] = 238;
assign img[ 8600] = 238;
assign img[ 8601] = 142;
assign img[ 8602] = 152;
assign img[ 8603] = 253;
assign img[ 8604] = 255;
assign img[ 8605] = 255;
assign img[ 8606] = 255;
assign img[ 8607] = 239;
assign img[ 8608] = 238;
assign img[ 8609] = 255;
assign img[ 8610] = 255;
assign img[ 8611] = 255;
assign img[ 8612] = 255;
assign img[ 8613] = 255;
assign img[ 8614] = 255;
assign img[ 8615] = 255;
assign img[ 8616] = 238;
assign img[ 8617] = 238;
assign img[ 8618] = 238;
assign img[ 8619] = 255;
assign img[ 8620] = 255;
assign img[ 8621] = 207;
assign img[ 8622] = 236;
assign img[ 8623] = 206;
assign img[ 8624] = 236;
assign img[ 8625] = 238;
assign img[ 8626] = 254;
assign img[ 8627] = 254;
assign img[ 8628] = 238;
assign img[ 8629] = 238;
assign img[ 8630] = 238;
assign img[ 8631] = 255;
assign img[ 8632] = 255;
assign img[ 8633] = 255;
assign img[ 8634] = 255;
assign img[ 8635] = 255;
assign img[ 8636] = 255;
assign img[ 8637] = 255;
assign img[ 8638] = 255;
assign img[ 8639] = 255;
assign img[ 8640] = 255;
assign img[ 8641] = 255;
assign img[ 8642] = 255;
assign img[ 8643] = 255;
assign img[ 8644] = 255;
assign img[ 8645] = 207;
assign img[ 8646] = 236;
assign img[ 8647] = 238;
assign img[ 8648] = 254;
assign img[ 8649] = 255;
assign img[ 8650] = 255;
assign img[ 8651] = 255;
assign img[ 8652] = 238;
assign img[ 8653] = 238;
assign img[ 8654] = 238;
assign img[ 8655] = 238;
assign img[ 8656] = 254;
assign img[ 8657] = 255;
assign img[ 8658] = 239;
assign img[ 8659] = 238;
assign img[ 8660] = 238;
assign img[ 8661] = 238;
assign img[ 8662] = 238;
assign img[ 8663] = 238;
assign img[ 8664] = 238;
assign img[ 8665] = 238;
assign img[ 8666] = 254;
assign img[ 8667] = 239;
assign img[ 8668] = 238;
assign img[ 8669] = 238;
assign img[ 8670] = 254;
assign img[ 8671] = 207;
assign img[ 8672] = 204;
assign img[ 8673] = 236;
assign img[ 8674] = 254;
assign img[ 8675] = 239;
assign img[ 8676] = 238;
assign img[ 8677] = 238;
assign img[ 8678] = 156;
assign img[ 8679] = 253;
assign img[ 8680] = 255;
assign img[ 8681] = 255;
assign img[ 8682] = 238;
assign img[ 8683] = 238;
assign img[ 8684] = 206;
assign img[ 8685] = 204;
assign img[ 8686] = 236;
assign img[ 8687] = 255;
assign img[ 8688] = 221;
assign img[ 8689] = 253;
assign img[ 8690] = 239;
assign img[ 8691] = 238;
assign img[ 8692] = 238;
assign img[ 8693] = 238;
assign img[ 8694] = 238;
assign img[ 8695] = 238;
assign img[ 8696] = 238;
assign img[ 8697] = 191;
assign img[ 8698] = 238;
assign img[ 8699] = 238;
assign img[ 8700] = 204;
assign img[ 8701] = 236;
assign img[ 8702] = 238;
assign img[ 8703] = 238;
assign img[ 8704] = 96;
assign img[ 8705] = 239;
assign img[ 8706] = 238;
assign img[ 8707] = 239;
assign img[ 8708] = 238;
assign img[ 8709] = 238;
assign img[ 8710] = 206;
assign img[ 8711] = 238;
assign img[ 8712] = 238;
assign img[ 8713] = 255;
assign img[ 8714] = 255;
assign img[ 8715] = 175;
assign img[ 8716] = 255;
assign img[ 8717] = 255;
assign img[ 8718] = 255;
assign img[ 8719] = 255;
assign img[ 8720] = 255;
assign img[ 8721] = 255;
assign img[ 8722] = 255;
assign img[ 8723] = 255;
assign img[ 8724] = 255;
assign img[ 8725] = 255;
assign img[ 8726] = 255;
assign img[ 8727] = 255;
assign img[ 8728] = 255;
assign img[ 8729] = 255;
assign img[ 8730] = 221;
assign img[ 8731] = 255;
assign img[ 8732] = 255;
assign img[ 8733] = 255;
assign img[ 8734] = 255;
assign img[ 8735] = 191;
assign img[ 8736] = 234;
assign img[ 8737] = 238;
assign img[ 8738] = 238;
assign img[ 8739] = 255;
assign img[ 8740] = 255;
assign img[ 8741] = 255;
assign img[ 8742] = 255;
assign img[ 8743] = 255;
assign img[ 8744] = 255;
assign img[ 8745] = 255;
assign img[ 8746] = 255;
assign img[ 8747] = 255;
assign img[ 8748] = 255;
assign img[ 8749] = 255;
assign img[ 8750] = 255;
assign img[ 8751] = 255;
assign img[ 8752] = 238;
assign img[ 8753] = 238;
assign img[ 8754] = 238;
assign img[ 8755] = 238;
assign img[ 8756] = 238;
assign img[ 8757] = 255;
assign img[ 8758] = 255;
assign img[ 8759] = 255;
assign img[ 8760] = 255;
assign img[ 8761] = 255;
assign img[ 8762] = 223;
assign img[ 8763] = 221;
assign img[ 8764] = 252;
assign img[ 8765] = 255;
assign img[ 8766] = 238;
assign img[ 8767] = 255;
assign img[ 8768] = 255;
assign img[ 8769] = 255;
assign img[ 8770] = 239;
assign img[ 8771] = 238;
assign img[ 8772] = 254;
assign img[ 8773] = 239;
assign img[ 8774] = 204;
assign img[ 8775] = 238;
assign img[ 8776] = 238;
assign img[ 8777] = 255;
assign img[ 8778] = 255;
assign img[ 8779] = 255;
assign img[ 8780] = 238;
assign img[ 8781] = 238;
assign img[ 8782] = 238;
assign img[ 8783] = 255;
assign img[ 8784] = 255;
assign img[ 8785] = 255;
assign img[ 8786] = 255;
assign img[ 8787] = 255;
assign img[ 8788] = 255;
assign img[ 8789] = 255;
assign img[ 8790] = 255;
assign img[ 8791] = 255;
assign img[ 8792] = 255;
assign img[ 8793] = 255;
assign img[ 8794] = 255;
assign img[ 8795] = 239;
assign img[ 8796] = 254;
assign img[ 8797] = 255;
assign img[ 8798] = 255;
assign img[ 8799] = 255;
assign img[ 8800] = 238;
assign img[ 8801] = 238;
assign img[ 8802] = 254;
assign img[ 8803] = 255;
assign img[ 8804] = 255;
assign img[ 8805] = 238;
assign img[ 8806] = 238;
assign img[ 8807] = 238;
assign img[ 8808] = 238;
assign img[ 8809] = 255;
assign img[ 8810] = 255;
assign img[ 8811] = 255;
assign img[ 8812] = 255;
assign img[ 8813] = 255;
assign img[ 8814] = 255;
assign img[ 8815] = 239;
assign img[ 8816] = 204;
assign img[ 8817] = 238;
assign img[ 8818] = 254;
assign img[ 8819] = 255;
assign img[ 8820] = 175;
assign img[ 8821] = 170;
assign img[ 8822] = 234;
assign img[ 8823] = 238;
assign img[ 8824] = 238;
assign img[ 8825] = 255;
assign img[ 8826] = 255;
assign img[ 8827] = 255;
assign img[ 8828] = 239;
assign img[ 8829] = 238;
assign img[ 8830] = 238;
assign img[ 8831] = 238;
assign img[ 8832] = 96;
assign img[ 8833] = 255;
assign img[ 8834] = 255;
assign img[ 8835] = 255;
assign img[ 8836] = 255;
assign img[ 8837] = 255;
assign img[ 8838] = 255;
assign img[ 8839] = 255;
assign img[ 8840] = 255;
assign img[ 8841] = 255;
assign img[ 8842] = 255;
assign img[ 8843] = 223;
assign img[ 8844] = 236;
assign img[ 8845] = 254;
assign img[ 8846] = 255;
assign img[ 8847] = 207;
assign img[ 8848] = 204;
assign img[ 8849] = 236;
assign img[ 8850] = 254;
assign img[ 8851] = 223;
assign img[ 8852] = 221;
assign img[ 8853] = 255;
assign img[ 8854] = 255;
assign img[ 8855] = 255;
assign img[ 8856] = 255;
assign img[ 8857] = 223;
assign img[ 8858] = 221;
assign img[ 8859] = 253;
assign img[ 8860] = 255;
assign img[ 8861] = 255;
assign img[ 8862] = 239;
assign img[ 8863] = 238;
assign img[ 8864] = 204;
assign img[ 8865] = 254;
assign img[ 8866] = 239;
assign img[ 8867] = 255;
assign img[ 8868] = 239;
assign img[ 8869] = 238;
assign img[ 8870] = 238;
assign img[ 8871] = 255;
assign img[ 8872] = 255;
assign img[ 8873] = 255;
assign img[ 8874] = 255;
assign img[ 8875] = 255;
assign img[ 8876] = 255;
assign img[ 8877] = 255;
assign img[ 8878] = 238;
assign img[ 8879] = 238;
assign img[ 8880] = 254;
assign img[ 8881] = 255;
assign img[ 8882] = 255;
assign img[ 8883] = 255;
assign img[ 8884] = 238;
assign img[ 8885] = 255;
assign img[ 8886] = 255;
assign img[ 8887] = 255;
assign img[ 8888] = 255;
assign img[ 8889] = 255;
assign img[ 8890] = 255;
assign img[ 8891] = 255;
assign img[ 8892] = 255;
assign img[ 8893] = 223;
assign img[ 8894] = 255;
assign img[ 8895] = 255;
assign img[ 8896] = 255;
assign img[ 8897] = 255;
assign img[ 8898] = 255;
assign img[ 8899] = 255;
assign img[ 8900] = 255;
assign img[ 8901] = 255;
assign img[ 8902] = 255;
assign img[ 8903] = 255;
assign img[ 8904] = 255;
assign img[ 8905] = 255;
assign img[ 8906] = 255;
assign img[ 8907] = 255;
assign img[ 8908] = 255;
assign img[ 8909] = 255;
assign img[ 8910] = 255;
assign img[ 8911] = 255;
assign img[ 8912] = 255;
assign img[ 8913] = 255;
assign img[ 8914] = 239;
assign img[ 8915] = 238;
assign img[ 8916] = 238;
assign img[ 8917] = 238;
assign img[ 8918] = 238;
assign img[ 8919] = 238;
assign img[ 8920] = 238;
assign img[ 8921] = 254;
assign img[ 8922] = 254;
assign img[ 8923] = 255;
assign img[ 8924] = 255;
assign img[ 8925] = 255;
assign img[ 8926] = 255;
assign img[ 8927] = 239;
assign img[ 8928] = 170;
assign img[ 8929] = 238;
assign img[ 8930] = 254;
assign img[ 8931] = 255;
assign img[ 8932] = 255;
assign img[ 8933] = 255;
assign img[ 8934] = 221;
assign img[ 8935] = 253;
assign img[ 8936] = 255;
assign img[ 8937] = 255;
assign img[ 8938] = 255;
assign img[ 8939] = 239;
assign img[ 8940] = 206;
assign img[ 8941] = 255;
assign img[ 8942] = 255;
assign img[ 8943] = 255;
assign img[ 8944] = 239;
assign img[ 8945] = 206;
assign img[ 8946] = 236;
assign img[ 8947] = 255;
assign img[ 8948] = 223;
assign img[ 8949] = 253;
assign img[ 8950] = 255;
assign img[ 8951] = 239;
assign img[ 8952] = 238;
assign img[ 8953] = 174;
assign img[ 8954] = 170;
assign img[ 8955] = 234;
assign img[ 8956] = 234;
assign img[ 8957] = 238;
assign img[ 8958] = 254;
assign img[ 8959] = 255;
assign img[ 8960] = 0;
assign img[ 8961] = 204;
assign img[ 8962] = 220;
assign img[ 8963] = 221;
assign img[ 8964] = 253;
assign img[ 8965] = 255;
assign img[ 8966] = 159;
assign img[ 8967] = 153;
assign img[ 8968] = 249;
assign img[ 8969] = 255;
assign img[ 8970] = 255;
assign img[ 8971] = 239;
assign img[ 8972] = 254;
assign img[ 8973] = 255;
assign img[ 8974] = 255;
assign img[ 8975] = 255;
assign img[ 8976] = 255;
assign img[ 8977] = 255;
assign img[ 8978] = 255;
assign img[ 8979] = 255;
assign img[ 8980] = 255;
assign img[ 8981] = 255;
assign img[ 8982] = 238;
assign img[ 8983] = 238;
assign img[ 8984] = 238;
assign img[ 8985] = 255;
assign img[ 8986] = 187;
assign img[ 8987] = 255;
assign img[ 8988] = 255;
assign img[ 8989] = 255;
assign img[ 8990] = 223;
assign img[ 8991] = 223;
assign img[ 8992] = 255;
assign img[ 8993] = 255;
assign img[ 8994] = 255;
assign img[ 8995] = 207;
assign img[ 8996] = 238;
assign img[ 8997] = 255;
assign img[ 8998] = 255;
assign img[ 8999] = 239;
assign img[ 9000] = 238;
assign img[ 9001] = 238;
assign img[ 9002] = 206;
assign img[ 9003] = 238;
assign img[ 9004] = 238;
assign img[ 9005] = 238;
assign img[ 9006] = 238;
assign img[ 9007] = 238;
assign img[ 9008] = 254;
assign img[ 9009] = 255;
assign img[ 9010] = 255;
assign img[ 9011] = 255;
assign img[ 9012] = 255;
assign img[ 9013] = 255;
assign img[ 9014] = 255;
assign img[ 9015] = 255;
assign img[ 9016] = 239;
assign img[ 9017] = 239;
assign img[ 9018] = 238;
assign img[ 9019] = 238;
assign img[ 9020] = 238;
assign img[ 9021] = 238;
assign img[ 9022] = 238;
assign img[ 9023] = 255;
assign img[ 9024] = 255;
assign img[ 9025] = 255;
assign img[ 9026] = 255;
assign img[ 9027] = 255;
assign img[ 9028] = 255;
assign img[ 9029] = 255;
assign img[ 9030] = 239;
assign img[ 9031] = 238;
assign img[ 9032] = 238;
assign img[ 9033] = 238;
assign img[ 9034] = 254;
assign img[ 9035] = 255;
assign img[ 9036] = 255;
assign img[ 9037] = 255;
assign img[ 9038] = 238;
assign img[ 9039] = 255;
assign img[ 9040] = 223;
assign img[ 9041] = 255;
assign img[ 9042] = 239;
assign img[ 9043] = 238;
assign img[ 9044] = 238;
assign img[ 9045] = 254;
assign img[ 9046] = 255;
assign img[ 9047] = 255;
assign img[ 9048] = 255;
assign img[ 9049] = 255;
assign img[ 9050] = 254;
assign img[ 9051] = 255;
assign img[ 9052] = 255;
assign img[ 9053] = 255;
assign img[ 9054] = 255;
assign img[ 9055] = 239;
assign img[ 9056] = 238;
assign img[ 9057] = 206;
assign img[ 9058] = 252;
assign img[ 9059] = 255;
assign img[ 9060] = 255;
assign img[ 9061] = 255;
assign img[ 9062] = 207;
assign img[ 9063] = 238;
assign img[ 9064] = 238;
assign img[ 9065] = 255;
assign img[ 9066] = 255;
assign img[ 9067] = 239;
assign img[ 9068] = 254;
assign img[ 9069] = 255;
assign img[ 9070] = 255;
assign img[ 9071] = 255;
assign img[ 9072] = 255;
assign img[ 9073] = 255;
assign img[ 9074] = 255;
assign img[ 9075] = 255;
assign img[ 9076] = 255;
assign img[ 9077] = 253;
assign img[ 9078] = 255;
assign img[ 9079] = 255;
assign img[ 9080] = 223;
assign img[ 9081] = 221;
assign img[ 9082] = 221;
assign img[ 9083] = 255;
assign img[ 9084] = 255;
assign img[ 9085] = 255;
assign img[ 9086] = 207;
assign img[ 9087] = 204;
assign img[ 9088] = 96;
assign img[ 9089] = 255;
assign img[ 9090] = 255;
assign img[ 9091] = 255;
assign img[ 9092] = 239;
assign img[ 9093] = 206;
assign img[ 9094] = 204;
assign img[ 9095] = 238;
assign img[ 9096] = 238;
assign img[ 9097] = 238;
assign img[ 9098] = 238;
assign img[ 9099] = 238;
assign img[ 9100] = 204;
assign img[ 9101] = 238;
assign img[ 9102] = 206;
assign img[ 9103] = 220;
assign img[ 9104] = 237;
assign img[ 9105] = 238;
assign img[ 9106] = 238;
assign img[ 9107] = 255;
assign img[ 9108] = 255;
assign img[ 9109] = 255;
assign img[ 9110] = 221;
assign img[ 9111] = 255;
assign img[ 9112] = 255;
assign img[ 9113] = 239;
assign img[ 9114] = 254;
assign img[ 9115] = 238;
assign img[ 9116] = 254;
assign img[ 9117] = 255;
assign img[ 9118] = 255;
assign img[ 9119] = 223;
assign img[ 9120] = 221;
assign img[ 9121] = 255;
assign img[ 9122] = 255;
assign img[ 9123] = 255;
assign img[ 9124] = 255;
assign img[ 9125] = 255;
assign img[ 9126] = 255;
assign img[ 9127] = 255;
assign img[ 9128] = 255;
assign img[ 9129] = 255;
assign img[ 9130] = 255;
assign img[ 9131] = 255;
assign img[ 9132] = 255;
assign img[ 9133] = 238;
assign img[ 9134] = 254;
assign img[ 9135] = 255;
assign img[ 9136] = 255;
assign img[ 9137] = 255;
assign img[ 9138] = 255;
assign img[ 9139] = 255;
assign img[ 9140] = 223;
assign img[ 9141] = 255;
assign img[ 9142] = 238;
assign img[ 9143] = 255;
assign img[ 9144] = 254;
assign img[ 9145] = 255;
assign img[ 9146] = 238;
assign img[ 9147] = 254;
assign img[ 9148] = 239;
assign img[ 9149] = 238;
assign img[ 9150] = 238;
assign img[ 9151] = 255;
assign img[ 9152] = 255;
assign img[ 9153] = 255;
assign img[ 9154] = 191;
assign img[ 9155] = 187;
assign img[ 9156] = 251;
assign img[ 9157] = 255;
assign img[ 9158] = 255;
assign img[ 9159] = 255;
assign img[ 9160] = 255;
assign img[ 9161] = 255;
assign img[ 9162] = 255;
assign img[ 9163] = 255;
assign img[ 9164] = 255;
assign img[ 9165] = 255;
assign img[ 9166] = 255;
assign img[ 9167] = 255;
assign img[ 9168] = 255;
assign img[ 9169] = 255;
assign img[ 9170] = 255;
assign img[ 9171] = 238;
assign img[ 9172] = 238;
assign img[ 9173] = 238;
assign img[ 9174] = 238;
assign img[ 9175] = 254;
assign img[ 9176] = 255;
assign img[ 9177] = 255;
assign img[ 9178] = 255;
assign img[ 9179] = 255;
assign img[ 9180] = 255;
assign img[ 9181] = 255;
assign img[ 9182] = 255;
assign img[ 9183] = 255;
assign img[ 9184] = 223;
assign img[ 9185] = 221;
assign img[ 9186] = 253;
assign img[ 9187] = 255;
assign img[ 9188] = 255;
assign img[ 9189] = 239;
assign img[ 9190] = 206;
assign img[ 9191] = 254;
assign img[ 9192] = 238;
assign img[ 9193] = 255;
assign img[ 9194] = 239;
assign img[ 9195] = 255;
assign img[ 9196] = 221;
assign img[ 9197] = 253;
assign img[ 9198] = 255;
assign img[ 9199] = 255;
assign img[ 9200] = 206;
assign img[ 9201] = 204;
assign img[ 9202] = 204;
assign img[ 9203] = 204;
assign img[ 9204] = 204;
assign img[ 9205] = 204;
assign img[ 9206] = 238;
assign img[ 9207] = 238;
assign img[ 9208] = 238;
assign img[ 9209] = 238;
assign img[ 9210] = 204;
assign img[ 9211] = 204;
assign img[ 9212] = 204;
assign img[ 9213] = 236;
assign img[ 9214] = 206;
assign img[ 9215] = 236;
assign img[ 9216] = 96;
assign img[ 9217] = 238;
assign img[ 9218] = 238;
assign img[ 9219] = 223;
assign img[ 9220] = 221;
assign img[ 9221] = 205;
assign img[ 9222] = 204;
assign img[ 9223] = 238;
assign img[ 9224] = 238;
assign img[ 9225] = 239;
assign img[ 9226] = 223;
assign img[ 9227] = 221;
assign img[ 9228] = 221;
assign img[ 9229] = 255;
assign img[ 9230] = 239;
assign img[ 9231] = 238;
assign img[ 9232] = 238;
assign img[ 9233] = 238;
assign img[ 9234] = 220;
assign img[ 9235] = 255;
assign img[ 9236] = 238;
assign img[ 9237] = 238;
assign img[ 9238] = 238;
assign img[ 9239] = 238;
assign img[ 9240] = 238;
assign img[ 9241] = 206;
assign img[ 9242] = 204;
assign img[ 9243] = 238;
assign img[ 9244] = 238;
assign img[ 9245] = 255;
assign img[ 9246] = 255;
assign img[ 9247] = 223;
assign img[ 9248] = 221;
assign img[ 9249] = 255;
assign img[ 9250] = 255;
assign img[ 9251] = 255;
assign img[ 9252] = 255;
assign img[ 9253] = 255;
assign img[ 9254] = 255;
assign img[ 9255] = 255;
assign img[ 9256] = 238;
assign img[ 9257] = 254;
assign img[ 9258] = 255;
assign img[ 9259] = 255;
assign img[ 9260] = 255;
assign img[ 9261] = 255;
assign img[ 9262] = 255;
assign img[ 9263] = 239;
assign img[ 9264] = 238;
assign img[ 9265] = 238;
assign img[ 9266] = 238;
assign img[ 9267] = 238;
assign img[ 9268] = 238;
assign img[ 9269] = 255;
assign img[ 9270] = 255;
assign img[ 9271] = 255;
assign img[ 9272] = 255;
assign img[ 9273] = 255;
assign img[ 9274] = 239;
assign img[ 9275] = 238;
assign img[ 9276] = 238;
assign img[ 9277] = 255;
assign img[ 9278] = 238;
assign img[ 9279] = 255;
assign img[ 9280] = 255;
assign img[ 9281] = 255;
assign img[ 9282] = 223;
assign img[ 9283] = 255;
assign img[ 9284] = 223;
assign img[ 9285] = 221;
assign img[ 9286] = 204;
assign img[ 9287] = 254;
assign img[ 9288] = 238;
assign img[ 9289] = 255;
assign img[ 9290] = 255;
assign img[ 9291] = 255;
assign img[ 9292] = 239;
assign img[ 9293] = 238;
assign img[ 9294] = 238;
assign img[ 9295] = 238;
assign img[ 9296] = 238;
assign img[ 9297] = 238;
assign img[ 9298] = 238;
assign img[ 9299] = 255;
assign img[ 9300] = 238;
assign img[ 9301] = 238;
assign img[ 9302] = 238;
assign img[ 9303] = 238;
assign img[ 9304] = 238;
assign img[ 9305] = 254;
assign img[ 9306] = 255;
assign img[ 9307] = 255;
assign img[ 9308] = 255;
assign img[ 9309] = 255;
assign img[ 9310] = 255;
assign img[ 9311] = 239;
assign img[ 9312] = 204;
assign img[ 9313] = 252;
assign img[ 9314] = 255;
assign img[ 9315] = 255;
assign img[ 9316] = 255;
assign img[ 9317] = 255;
assign img[ 9318] = 255;
assign img[ 9319] = 255;
assign img[ 9320] = 255;
assign img[ 9321] = 239;
assign img[ 9322] = 238;
assign img[ 9323] = 239;
assign img[ 9324] = 238;
assign img[ 9325] = 238;
assign img[ 9326] = 206;
assign img[ 9327] = 238;
assign img[ 9328] = 238;
assign img[ 9329] = 239;
assign img[ 9330] = 255;
assign img[ 9331] = 239;
assign img[ 9332] = 254;
assign img[ 9333] = 223;
assign img[ 9334] = 237;
assign img[ 9335] = 238;
assign img[ 9336] = 238;
assign img[ 9337] = 174;
assign img[ 9338] = 170;
assign img[ 9339] = 255;
assign img[ 9340] = 238;
assign img[ 9341] = 238;
assign img[ 9342] = 254;
assign img[ 9343] = 255;
assign img[ 9344] = 96;
assign img[ 9345] = 223;
assign img[ 9346] = 253;
assign img[ 9347] = 239;
assign img[ 9348] = 238;
assign img[ 9349] = 238;
assign img[ 9350] = 238;
assign img[ 9351] = 255;
assign img[ 9352] = 255;
assign img[ 9353] = 255;
assign img[ 9354] = 255;
assign img[ 9355] = 255;
assign img[ 9356] = 221;
assign img[ 9357] = 253;
assign img[ 9358] = 238;
assign img[ 9359] = 255;
assign img[ 9360] = 255;
assign img[ 9361] = 255;
assign img[ 9362] = 255;
assign img[ 9363] = 255;
assign img[ 9364] = 221;
assign img[ 9365] = 253;
assign img[ 9366] = 255;
assign img[ 9367] = 255;
assign img[ 9368] = 255;
assign img[ 9369] = 255;
assign img[ 9370] = 187;
assign img[ 9371] = 171;
assign img[ 9372] = 234;
assign img[ 9373] = 238;
assign img[ 9374] = 206;
assign img[ 9375] = 174;
assign img[ 9376] = 170;
assign img[ 9377] = 238;
assign img[ 9378] = 238;
assign img[ 9379] = 255;
assign img[ 9380] = 238;
assign img[ 9381] = 238;
assign img[ 9382] = 238;
assign img[ 9383] = 255;
assign img[ 9384] = 255;
assign img[ 9385] = 255;
assign img[ 9386] = 221;
assign img[ 9387] = 255;
assign img[ 9388] = 255;
assign img[ 9389] = 239;
assign img[ 9390] = 238;
assign img[ 9391] = 238;
assign img[ 9392] = 238;
assign img[ 9393] = 238;
assign img[ 9394] = 254;
assign img[ 9395] = 255;
assign img[ 9396] = 255;
assign img[ 9397] = 255;
assign img[ 9398] = 255;
assign img[ 9399] = 255;
assign img[ 9400] = 255;
assign img[ 9401] = 255;
assign img[ 9402] = 221;
assign img[ 9403] = 253;
assign img[ 9404] = 254;
assign img[ 9405] = 255;
assign img[ 9406] = 254;
assign img[ 9407] = 255;
assign img[ 9408] = 254;
assign img[ 9409] = 255;
assign img[ 9410] = 255;
assign img[ 9411] = 255;
assign img[ 9412] = 255;
assign img[ 9413] = 255;
assign img[ 9414] = 255;
assign img[ 9415] = 255;
assign img[ 9416] = 255;
assign img[ 9417] = 255;
assign img[ 9418] = 255;
assign img[ 9419] = 255;
assign img[ 9420] = 255;
assign img[ 9421] = 255;
assign img[ 9422] = 255;
assign img[ 9423] = 255;
assign img[ 9424] = 255;
assign img[ 9425] = 255;
assign img[ 9426] = 255;
assign img[ 9427] = 255;
assign img[ 9428] = 255;
assign img[ 9429] = 255;
assign img[ 9430] = 255;
assign img[ 9431] = 255;
assign img[ 9432] = 255;
assign img[ 9433] = 239;
assign img[ 9434] = 238;
assign img[ 9435] = 238;
assign img[ 9436] = 238;
assign img[ 9437] = 238;
assign img[ 9438] = 238;
assign img[ 9439] = 238;
assign img[ 9440] = 254;
assign img[ 9441] = 223;
assign img[ 9442] = 253;
assign img[ 9443] = 223;
assign img[ 9444] = 221;
assign img[ 9445] = 221;
assign img[ 9446] = 189;
assign img[ 9447] = 255;
assign img[ 9448] = 255;
assign img[ 9449] = 255;
assign img[ 9450] = 255;
assign img[ 9451] = 255;
assign img[ 9452] = 221;
assign img[ 9453] = 253;
assign img[ 9454] = 255;
assign img[ 9455] = 191;
assign img[ 9456] = 187;
assign img[ 9457] = 255;
assign img[ 9458] = 255;
assign img[ 9459] = 255;
assign img[ 9460] = 221;
assign img[ 9461] = 237;
assign img[ 9462] = 238;
assign img[ 9463] = 238;
assign img[ 9464] = 238;
assign img[ 9465] = 255;
assign img[ 9466] = 255;
assign img[ 9467] = 255;
assign img[ 9468] = 223;
assign img[ 9469] = 255;
assign img[ 9470] = 255;
assign img[ 9471] = 255;
assign img[ 9472] = 96;
assign img[ 9473] = 238;
assign img[ 9474] = 254;
assign img[ 9475] = 239;
assign img[ 9476] = 204;
assign img[ 9477] = 204;
assign img[ 9478] = 204;
assign img[ 9479] = 220;
assign img[ 9480] = 253;
assign img[ 9481] = 255;
assign img[ 9482] = 238;
assign img[ 9483] = 255;
assign img[ 9484] = 255;
assign img[ 9485] = 255;
assign img[ 9486] = 255;
assign img[ 9487] = 223;
assign img[ 9488] = 253;
assign img[ 9489] = 255;
assign img[ 9490] = 255;
assign img[ 9491] = 207;
assign img[ 9492] = 220;
assign img[ 9493] = 253;
assign img[ 9494] = 255;
assign img[ 9495] = 255;
assign img[ 9496] = 255;
assign img[ 9497] = 255;
assign img[ 9498] = 255;
assign img[ 9499] = 223;
assign img[ 9500] = 253;
assign img[ 9501] = 255;
assign img[ 9502] = 255;
assign img[ 9503] = 255;
assign img[ 9504] = 255;
assign img[ 9505] = 255;
assign img[ 9506] = 239;
assign img[ 9507] = 238;
assign img[ 9508] = 238;
assign img[ 9509] = 238;
assign img[ 9510] = 238;
assign img[ 9511] = 255;
assign img[ 9512] = 255;
assign img[ 9513] = 255;
assign img[ 9514] = 191;
assign img[ 9515] = 255;
assign img[ 9516] = 255;
assign img[ 9517] = 255;
assign img[ 9518] = 255;
assign img[ 9519] = 255;
assign img[ 9520] = 255;
assign img[ 9521] = 255;
assign img[ 9522] = 255;
assign img[ 9523] = 255;
assign img[ 9524] = 205;
assign img[ 9525] = 238;
assign img[ 9526] = 238;
assign img[ 9527] = 238;
assign img[ 9528] = 238;
assign img[ 9529] = 238;
assign img[ 9530] = 206;
assign img[ 9531] = 221;
assign img[ 9532] = 236;
assign img[ 9533] = 238;
assign img[ 9534] = 238;
assign img[ 9535] = 254;
assign img[ 9536] = 255;
assign img[ 9537] = 191;
assign img[ 9538] = 187;
assign img[ 9539] = 255;
assign img[ 9540] = 239;
assign img[ 9541] = 238;
assign img[ 9542] = 238;
assign img[ 9543] = 254;
assign img[ 9544] = 255;
assign img[ 9545] = 255;
assign img[ 9546] = 238;
assign img[ 9547] = 255;
assign img[ 9548] = 255;
assign img[ 9549] = 255;
assign img[ 9550] = 255;
assign img[ 9551] = 255;
assign img[ 9552] = 255;
assign img[ 9553] = 255;
assign img[ 9554] = 255;
assign img[ 9555] = 255;
assign img[ 9556] = 255;
assign img[ 9557] = 255;
assign img[ 9558] = 255;
assign img[ 9559] = 255;
assign img[ 9560] = 255;
assign img[ 9561] = 255;
assign img[ 9562] = 255;
assign img[ 9563] = 255;
assign img[ 9564] = 254;
assign img[ 9565] = 255;
assign img[ 9566] = 238;
assign img[ 9567] = 206;
assign img[ 9568] = 236;
assign img[ 9569] = 254;
assign img[ 9570] = 255;
assign img[ 9571] = 255;
assign img[ 9572] = 223;
assign img[ 9573] = 221;
assign img[ 9574] = 253;
assign img[ 9575] = 255;
assign img[ 9576] = 255;
assign img[ 9577] = 255;
assign img[ 9578] = 238;
assign img[ 9579] = 255;
assign img[ 9580] = 221;
assign img[ 9581] = 253;
assign img[ 9582] = 223;
assign img[ 9583] = 253;
assign img[ 9584] = 223;
assign img[ 9585] = 253;
assign img[ 9586] = 255;
assign img[ 9587] = 255;
assign img[ 9588] = 205;
assign img[ 9589] = 238;
assign img[ 9590] = 254;
assign img[ 9591] = 255;
assign img[ 9592] = 255;
assign img[ 9593] = 191;
assign img[ 9594] = 187;
assign img[ 9595] = 155;
assign img[ 9596] = 217;
assign img[ 9597] = 253;
assign img[ 9598] = 255;
assign img[ 9599] = 255;
assign img[ 9600] = 64;
assign img[ 9601] = 204;
assign img[ 9602] = 236;
assign img[ 9603] = 206;
assign img[ 9604] = 236;
assign img[ 9605] = 254;
assign img[ 9606] = 255;
assign img[ 9607] = 239;
assign img[ 9608] = 238;
assign img[ 9609] = 238;
assign img[ 9610] = 206;
assign img[ 9611] = 205;
assign img[ 9612] = 236;
assign img[ 9613] = 238;
assign img[ 9614] = 238;
assign img[ 9615] = 206;
assign img[ 9616] = 204;
assign img[ 9617] = 238;
assign img[ 9618] = 238;
assign img[ 9619] = 254;
assign img[ 9620] = 238;
assign img[ 9621] = 255;
assign img[ 9622] = 238;
assign img[ 9623] = 254;
assign img[ 9624] = 255;
assign img[ 9625] = 255;
assign img[ 9626] = 170;
assign img[ 9627] = 251;
assign img[ 9628] = 239;
assign img[ 9629] = 255;
assign img[ 9630] = 255;
assign img[ 9631] = 191;
assign img[ 9632] = 187;
assign img[ 9633] = 255;
assign img[ 9634] = 255;
assign img[ 9635] = 255;
assign img[ 9636] = 191;
assign img[ 9637] = 171;
assign img[ 9638] = 234;
assign img[ 9639] = 255;
assign img[ 9640] = 255;
assign img[ 9641] = 255;
assign img[ 9642] = 255;
assign img[ 9643] = 255;
assign img[ 9644] = 255;
assign img[ 9645] = 238;
assign img[ 9646] = 238;
assign img[ 9647] = 254;
assign img[ 9648] = 238;
assign img[ 9649] = 255;
assign img[ 9650] = 254;
assign img[ 9651] = 255;
assign img[ 9652] = 255;
assign img[ 9653] = 255;
assign img[ 9654] = 255;
assign img[ 9655] = 255;
assign img[ 9656] = 255;
assign img[ 9657] = 255;
assign img[ 9658] = 239;
assign img[ 9659] = 254;
assign img[ 9660] = 255;
assign img[ 9661] = 255;
assign img[ 9662] = 255;
assign img[ 9663] = 255;
assign img[ 9664] = 255;
assign img[ 9665] = 255;
assign img[ 9666] = 255;
assign img[ 9667] = 255;
assign img[ 9668] = 255;
assign img[ 9669] = 255;
assign img[ 9670] = 255;
assign img[ 9671] = 255;
assign img[ 9672] = 255;
assign img[ 9673] = 255;
assign img[ 9674] = 255;
assign img[ 9675] = 255;
assign img[ 9676] = 239;
assign img[ 9677] = 238;
assign img[ 9678] = 238;
assign img[ 9679] = 238;
assign img[ 9680] = 238;
assign img[ 9681] = 254;
assign img[ 9682] = 238;
assign img[ 9683] = 238;
assign img[ 9684] = 204;
assign img[ 9685] = 204;
assign img[ 9686] = 238;
assign img[ 9687] = 238;
assign img[ 9688] = 238;
assign img[ 9689] = 254;
assign img[ 9690] = 238;
assign img[ 9691] = 174;
assign img[ 9692] = 250;
assign img[ 9693] = 255;
assign img[ 9694] = 255;
assign img[ 9695] = 206;
assign img[ 9696] = 140;
assign img[ 9697] = 170;
assign img[ 9698] = 250;
assign img[ 9699] = 255;
assign img[ 9700] = 238;
assign img[ 9701] = 255;
assign img[ 9702] = 255;
assign img[ 9703] = 255;
assign img[ 9704] = 255;
assign img[ 9705] = 255;
assign img[ 9706] = 238;
assign img[ 9707] = 254;
assign img[ 9708] = 255;
assign img[ 9709] = 255;
assign img[ 9710] = 255;
assign img[ 9711] = 255;
assign img[ 9712] = 255;
assign img[ 9713] = 255;
assign img[ 9714] = 255;
assign img[ 9715] = 239;
assign img[ 9716] = 206;
assign img[ 9717] = 220;
assign img[ 9718] = 253;
assign img[ 9719] = 255;
assign img[ 9720] = 255;
assign img[ 9721] = 255;
assign img[ 9722] = 187;
assign img[ 9723] = 255;
assign img[ 9724] = 255;
assign img[ 9725] = 255;
assign img[ 9726] = 223;
assign img[ 9727] = 221;
assign img[ 9728] = 32;
assign img[ 9729] = 238;
assign img[ 9730] = 238;
assign img[ 9731] = 255;
assign img[ 9732] = 141;
assign img[ 9733] = 170;
assign img[ 9734] = 250;
assign img[ 9735] = 255;
assign img[ 9736] = 255;
assign img[ 9737] = 255;
assign img[ 9738] = 238;
assign img[ 9739] = 238;
assign img[ 9740] = 222;
assign img[ 9741] = 255;
assign img[ 9742] = 255;
assign img[ 9743] = 255;
assign img[ 9744] = 187;
assign img[ 9745] = 255;
assign img[ 9746] = 253;
assign img[ 9747] = 253;
assign img[ 9748] = 238;
assign img[ 9749] = 254;
assign img[ 9750] = 238;
assign img[ 9751] = 238;
assign img[ 9752] = 238;
assign img[ 9753] = 207;
assign img[ 9754] = 204;
assign img[ 9755] = 236;
assign img[ 9756] = 238;
assign img[ 9757] = 255;
assign img[ 9758] = 255;
assign img[ 9759] = 255;
assign img[ 9760] = 155;
assign img[ 9761] = 255;
assign img[ 9762] = 255;
assign img[ 9763] = 255;
assign img[ 9764] = 223;
assign img[ 9765] = 255;
assign img[ 9766] = 255;
assign img[ 9767] = 255;
assign img[ 9768] = 238;
assign img[ 9769] = 238;
assign img[ 9770] = 238;
assign img[ 9771] = 238;
assign img[ 9772] = 238;
assign img[ 9773] = 206;
assign img[ 9774] = 236;
assign img[ 9775] = 223;
assign img[ 9776] = 253;
assign img[ 9777] = 255;
assign img[ 9778] = 255;
assign img[ 9779] = 255;
assign img[ 9780] = 239;
assign img[ 9781] = 254;
assign img[ 9782] = 255;
assign img[ 9783] = 255;
assign img[ 9784] = 255;
assign img[ 9785] = 255;
assign img[ 9786] = 255;
assign img[ 9787] = 255;
assign img[ 9788] = 238;
assign img[ 9789] = 255;
assign img[ 9790] = 254;
assign img[ 9791] = 255;
assign img[ 9792] = 255;
assign img[ 9793] = 255;
assign img[ 9794] = 191;
assign img[ 9795] = 255;
assign img[ 9796] = 255;
assign img[ 9797] = 255;
assign img[ 9798] = 223;
assign img[ 9799] = 255;
assign img[ 9800] = 255;
assign img[ 9801] = 239;
assign img[ 9802] = 254;
assign img[ 9803] = 255;
assign img[ 9804] = 238;
assign img[ 9805] = 238;
assign img[ 9806] = 238;
assign img[ 9807] = 255;
assign img[ 9808] = 207;
assign img[ 9809] = 238;
assign img[ 9810] = 222;
assign img[ 9811] = 221;
assign img[ 9812] = 236;
assign img[ 9813] = 238;
assign img[ 9814] = 238;
assign img[ 9815] = 254;
assign img[ 9816] = 255;
assign img[ 9817] = 255;
assign img[ 9818] = 254;
assign img[ 9819] = 206;
assign img[ 9820] = 254;
assign img[ 9821] = 255;
assign img[ 9822] = 255;
assign img[ 9823] = 255;
assign img[ 9824] = 255;
assign img[ 9825] = 255;
assign img[ 9826] = 255;
assign img[ 9827] = 255;
assign img[ 9828] = 255;
assign img[ 9829] = 207;
assign img[ 9830] = 238;
assign img[ 9831] = 238;
assign img[ 9832] = 238;
assign img[ 9833] = 255;
assign img[ 9834] = 255;
assign img[ 9835] = 255;
assign img[ 9836] = 239;
assign img[ 9837] = 254;
assign img[ 9838] = 255;
assign img[ 9839] = 255;
assign img[ 9840] = 255;
assign img[ 9841] = 255;
assign img[ 9842] = 255;
assign img[ 9843] = 223;
assign img[ 9844] = 221;
assign img[ 9845] = 221;
assign img[ 9846] = 236;
assign img[ 9847] = 254;
assign img[ 9848] = 254;
assign img[ 9849] = 223;
assign img[ 9850] = 221;
assign img[ 9851] = 221;
assign img[ 9852] = 153;
assign img[ 9853] = 255;
assign img[ 9854] = 255;
assign img[ 9855] = 255;
assign img[ 9856] = 96;
assign img[ 9857] = 239;
assign img[ 9858] = 255;
assign img[ 9859] = 223;
assign img[ 9860] = 221;
assign img[ 9861] = 255;
assign img[ 9862] = 223;
assign img[ 9863] = 255;
assign img[ 9864] = 255;
assign img[ 9865] = 255;
assign img[ 9866] = 239;
assign img[ 9867] = 238;
assign img[ 9868] = 238;
assign img[ 9869] = 238;
assign img[ 9870] = 238;
assign img[ 9871] = 254;
assign img[ 9872] = 220;
assign img[ 9873] = 255;
assign img[ 9874] = 255;
assign img[ 9875] = 239;
assign img[ 9876] = 238;
assign img[ 9877] = 238;
assign img[ 9878] = 238;
assign img[ 9879] = 238;
assign img[ 9880] = 254;
assign img[ 9881] = 239;
assign img[ 9882] = 170;
assign img[ 9883] = 238;
assign img[ 9884] = 238;
assign img[ 9885] = 255;
assign img[ 9886] = 223;
assign img[ 9887] = 221;
assign img[ 9888] = 221;
assign img[ 9889] = 253;
assign img[ 9890] = 255;
assign img[ 9891] = 255;
assign img[ 9892] = 255;
assign img[ 9893] = 255;
assign img[ 9894] = 255;
assign img[ 9895] = 255;
assign img[ 9896] = 238;
assign img[ 9897] = 238;
assign img[ 9898] = 206;
assign img[ 9899] = 255;
assign img[ 9900] = 255;
assign img[ 9901] = 255;
assign img[ 9902] = 238;
assign img[ 9903] = 238;
assign img[ 9904] = 254;
assign img[ 9905] = 255;
assign img[ 9906] = 255;
assign img[ 9907] = 255;
assign img[ 9908] = 223;
assign img[ 9909] = 255;
assign img[ 9910] = 255;
assign img[ 9911] = 255;
assign img[ 9912] = 207;
assign img[ 9913] = 204;
assign img[ 9914] = 204;
assign img[ 9915] = 238;
assign img[ 9916] = 254;
assign img[ 9917] = 239;
assign img[ 9918] = 238;
assign img[ 9919] = 255;
assign img[ 9920] = 255;
assign img[ 9921] = 255;
assign img[ 9922] = 255;
assign img[ 9923] = 255;
assign img[ 9924] = 255;
assign img[ 9925] = 239;
assign img[ 9926] = 254;
assign img[ 9927] = 223;
assign img[ 9928] = 238;
assign img[ 9929] = 238;
assign img[ 9930] = 255;
assign img[ 9931] = 223;
assign img[ 9932] = 221;
assign img[ 9933] = 255;
assign img[ 9934] = 255;
assign img[ 9935] = 255;
assign img[ 9936] = 255;
assign img[ 9937] = 255;
assign img[ 9938] = 239;
assign img[ 9939] = 238;
assign img[ 9940] = 238;
assign img[ 9941] = 255;
assign img[ 9942] = 255;
assign img[ 9943] = 255;
assign img[ 9944] = 239;
assign img[ 9945] = 254;
assign img[ 9946] = 255;
assign img[ 9947] = 255;
assign img[ 9948] = 255;
assign img[ 9949] = 255;
assign img[ 9950] = 255;
assign img[ 9951] = 255;
assign img[ 9952] = 255;
assign img[ 9953] = 255;
assign img[ 9954] = 255;
assign img[ 9955] = 255;
assign img[ 9956] = 255;
assign img[ 9957] = 239;
assign img[ 9958] = 238;
assign img[ 9959] = 238;
assign img[ 9960] = 238;
assign img[ 9961] = 255;
assign img[ 9962] = 238;
assign img[ 9963] = 255;
assign img[ 9964] = 238;
assign img[ 9965] = 238;
assign img[ 9966] = 238;
assign img[ 9967] = 255;
assign img[ 9968] = 255;
assign img[ 9969] = 255;
assign img[ 9970] = 238;
assign img[ 9971] = 255;
assign img[ 9972] = 238;
assign img[ 9973] = 238;
assign img[ 9974] = 238;
assign img[ 9975] = 238;
assign img[ 9976] = 238;
assign img[ 9977] = 238;
assign img[ 9978] = 204;
assign img[ 9979] = 204;
assign img[ 9980] = 238;
assign img[ 9981] = 255;
assign img[ 9982] = 207;
assign img[ 9983] = 236;
assign img[ 9984] = 0;
assign img[ 9985] = 198;
assign img[ 9986] = 238;
assign img[ 9987] = 255;
assign img[ 9988] = 153;
assign img[ 9989] = 153;
assign img[ 9990] = 185;
assign img[ 9991] = 155;
assign img[ 9992] = 249;
assign img[ 9993] = 255;
assign img[ 9994] = 255;
assign img[ 9995] = 255;
assign img[ 9996] = 238;
assign img[ 9997] = 238;
assign img[ 9998] = 254;
assign img[ 9999] = 255;
assign img[10000] = 255;
assign img[10001] = 255;
assign img[10002] = 255;
assign img[10003] = 255;
assign img[10004] = 223;
assign img[10005] = 255;
assign img[10006] = 255;
assign img[10007] = 255;
assign img[10008] = 255;
assign img[10009] = 255;
assign img[10010] = 255;
assign img[10011] = 255;
assign img[10012] = 255;
assign img[10013] = 255;
assign img[10014] = 255;
assign img[10015] = 223;
assign img[10016] = 255;
assign img[10017] = 255;
assign img[10018] = 255;
assign img[10019] = 255;
assign img[10020] = 255;
assign img[10021] = 255;
assign img[10022] = 255;
assign img[10023] = 255;
assign img[10024] = 238;
assign img[10025] = 238;
assign img[10026] = 238;
assign img[10027] = 238;
assign img[10028] = 170;
assign img[10029] = 250;
assign img[10030] = 255;
assign img[10031] = 255;
assign img[10032] = 255;
assign img[10033] = 255;
assign img[10034] = 255;
assign img[10035] = 255;
assign img[10036] = 255;
assign img[10037] = 255;
assign img[10038] = 255;
assign img[10039] = 255;
assign img[10040] = 255;
assign img[10041] = 239;
assign img[10042] = 206;
assign img[10043] = 238;
assign img[10044] = 238;
assign img[10045] = 255;
assign img[10046] = 255;
assign img[10047] = 255;
assign img[10048] = 255;
assign img[10049] = 255;
assign img[10050] = 223;
assign img[10051] = 255;
assign img[10052] = 255;
assign img[10053] = 223;
assign img[10054] = 221;
assign img[10055] = 254;
assign img[10056] = 254;
assign img[10057] = 255;
assign img[10058] = 255;
assign img[10059] = 255;
assign img[10060] = 255;
assign img[10061] = 255;
assign img[10062] = 255;
assign img[10063] = 255;
assign img[10064] = 255;
assign img[10065] = 255;
assign img[10066] = 255;
assign img[10067] = 239;
assign img[10068] = 254;
assign img[10069] = 255;
assign img[10070] = 238;
assign img[10071] = 238;
assign img[10072] = 238;
assign img[10073] = 255;
assign img[10074] = 223;
assign img[10075] = 255;
assign img[10076] = 255;
assign img[10077] = 255;
assign img[10078] = 255;
assign img[10079] = 255;
assign img[10080] = 204;
assign img[10081] = 204;
assign img[10082] = 253;
assign img[10083] = 255;
assign img[10084] = 255;
assign img[10085] = 255;
assign img[10086] = 255;
assign img[10087] = 255;
assign img[10088] = 255;
assign img[10089] = 255;
assign img[10090] = 255;
assign img[10091] = 239;
assign img[10092] = 220;
assign img[10093] = 255;
assign img[10094] = 255;
assign img[10095] = 255;
assign img[10096] = 221;
assign img[10097] = 221;
assign img[10098] = 253;
assign img[10099] = 255;
assign img[10100] = 239;
assign img[10101] = 238;
assign img[10102] = 238;
assign img[10103] = 238;
assign img[10104] = 238;
assign img[10105] = 174;
assign img[10106] = 138;
assign img[10107] = 136;
assign img[10108] = 136;
assign img[10109] = 234;
assign img[10110] = 238;
assign img[10111] = 254;
assign img[10112] = 96;
assign img[10113] = 239;
assign img[10114] = 238;
assign img[10115] = 255;
assign img[10116] = 238;
assign img[10117] = 238;
assign img[10118] = 206;
assign img[10119] = 204;
assign img[10120] = 236;
assign img[10121] = 238;
assign img[10122] = 206;
assign img[10123] = 204;
assign img[10124] = 236;
assign img[10125] = 238;
assign img[10126] = 238;
assign img[10127] = 255;
assign img[10128] = 255;
assign img[10129] = 255;
assign img[10130] = 255;
assign img[10131] = 255;
assign img[10132] = 239;
assign img[10133] = 238;
assign img[10134] = 254;
assign img[10135] = 255;
assign img[10136] = 255;
assign img[10137] = 175;
assign img[10138] = 138;
assign img[10139] = 238;
assign img[10140] = 238;
assign img[10141] = 255;
assign img[10142] = 255;
assign img[10143] = 239;
assign img[10144] = 238;
assign img[10145] = 238;
assign img[10146] = 238;
assign img[10147] = 255;
assign img[10148] = 255;
assign img[10149] = 255;
assign img[10150] = 255;
assign img[10151] = 255;
assign img[10152] = 255;
assign img[10153] = 255;
assign img[10154] = 255;
assign img[10155] = 207;
assign img[10156] = 236;
assign img[10157] = 238;
assign img[10158] = 238;
assign img[10159] = 239;
assign img[10160] = 255;
assign img[10161] = 255;
assign img[10162] = 255;
assign img[10163] = 255;
assign img[10164] = 255;
assign img[10165] = 255;
assign img[10166] = 255;
assign img[10167] = 255;
assign img[10168] = 255;
assign img[10169] = 255;
assign img[10170] = 223;
assign img[10171] = 255;
assign img[10172] = 255;
assign img[10173] = 255;
assign img[10174] = 255;
assign img[10175] = 255;
assign img[10176] = 255;
assign img[10177] = 239;
assign img[10178] = 238;
assign img[10179] = 238;
assign img[10180] = 254;
assign img[10181] = 255;
assign img[10182] = 255;
assign img[10183] = 255;
assign img[10184] = 255;
assign img[10185] = 255;
assign img[10186] = 255;
assign img[10187] = 255;
assign img[10188] = 255;
assign img[10189] = 255;
assign img[10190] = 255;
assign img[10191] = 255;
assign img[10192] = 255;
assign img[10193] = 255;
assign img[10194] = 223;
assign img[10195] = 255;
assign img[10196] = 255;
assign img[10197] = 223;
assign img[10198] = 253;
assign img[10199] = 255;
assign img[10200] = 255;
assign img[10201] = 255;
assign img[10202] = 255;
assign img[10203] = 255;
assign img[10204] = 255;
assign img[10205] = 255;
assign img[10206] = 255;
assign img[10207] = 239;
assign img[10208] = 238;
assign img[10209] = 238;
assign img[10210] = 254;
assign img[10211] = 255;
assign img[10212] = 255;
assign img[10213] = 238;
assign img[10214] = 204;
assign img[10215] = 238;
assign img[10216] = 254;
assign img[10217] = 239;
assign img[10218] = 238;
assign img[10219] = 238;
assign img[10220] = 255;
assign img[10221] = 255;
assign img[10222] = 255;
assign img[10223] = 255;
assign img[10224] = 255;
assign img[10225] = 255;
assign img[10226] = 255;
assign img[10227] = 255;
assign img[10228] = 223;
assign img[10229] = 221;
assign img[10230] = 236;
assign img[10231] = 254;
assign img[10232] = 255;
assign img[10233] = 255;
assign img[10234] = 236;
assign img[10235] = 223;
assign img[10236] = 204;
assign img[10237] = 238;
assign img[10238] = 238;
assign img[10239] = 238;
assign img[10240] = 96;
assign img[10241] = 206;
assign img[10242] = 252;
assign img[10243] = 223;
assign img[10244] = 189;
assign img[10245] = 171;
assign img[10246] = 170;
assign img[10247] = 234;
assign img[10248] = 238;
assign img[10249] = 238;
assign img[10250] = 238;
assign img[10251] = 238;
assign img[10252] = 254;
assign img[10253] = 255;
assign img[10254] = 255;
assign img[10255] = 255;
assign img[10256] = 238;
assign img[10257] = 255;
assign img[10258] = 255;
assign img[10259] = 255;
assign img[10260] = 238;
assign img[10261] = 238;
assign img[10262] = 238;
assign img[10263] = 254;
assign img[10264] = 255;
assign img[10265] = 255;
assign img[10266] = 238;
assign img[10267] = 238;
assign img[10268] = 238;
assign img[10269] = 255;
assign img[10270] = 255;
assign img[10271] = 191;
assign img[10272] = 238;
assign img[10273] = 254;
assign img[10274] = 255;
assign img[10275] = 255;
assign img[10276] = 255;
assign img[10277] = 255;
assign img[10278] = 255;
assign img[10279] = 255;
assign img[10280] = 255;
assign img[10281] = 255;
assign img[10282] = 223;
assign img[10283] = 221;
assign img[10284] = 253;
assign img[10285] = 239;
assign img[10286] = 238;
assign img[10287] = 238;
assign img[10288] = 254;
assign img[10289] = 255;
assign img[10290] = 221;
assign img[10291] = 253;
assign img[10292] = 255;
assign img[10293] = 255;
assign img[10294] = 255;
assign img[10295] = 255;
assign img[10296] = 255;
assign img[10297] = 255;
assign img[10298] = 206;
assign img[10299] = 255;
assign img[10300] = 255;
assign img[10301] = 255;
assign img[10302] = 238;
assign img[10303] = 238;
assign img[10304] = 238;
assign img[10305] = 239;
assign img[10306] = 238;
assign img[10307] = 238;
assign img[10308] = 254;
assign img[10309] = 255;
assign img[10310] = 255;
assign img[10311] = 255;
assign img[10312] = 255;
assign img[10313] = 255;
assign img[10314] = 255;
assign img[10315] = 239;
assign img[10316] = 254;
assign img[10317] = 223;
assign img[10318] = 221;
assign img[10319] = 255;
assign img[10320] = 255;
assign img[10321] = 255;
assign img[10322] = 255;
assign img[10323] = 255;
assign img[10324] = 255;
assign img[10325] = 207;
assign img[10326] = 236;
assign img[10327] = 238;
assign img[10328] = 222;
assign img[10329] = 221;
assign img[10330] = 253;
assign img[10331] = 255;
assign img[10332] = 255;
assign img[10333] = 255;
assign img[10334] = 255;
assign img[10335] = 255;
assign img[10336] = 238;
assign img[10337] = 238;
assign img[10338] = 254;
assign img[10339] = 255;
assign img[10340] = 223;
assign img[10341] = 255;
assign img[10342] = 255;
assign img[10343] = 255;
assign img[10344] = 255;
assign img[10345] = 255;
assign img[10346] = 255;
assign img[10347] = 239;
assign img[10348] = 206;
assign img[10349] = 238;
assign img[10350] = 238;
assign img[10351] = 255;
assign img[10352] = 239;
assign img[10353] = 238;
assign img[10354] = 238;
assign img[10355] = 238;
assign img[10356] = 204;
assign img[10357] = 238;
assign img[10358] = 238;
assign img[10359] = 255;
assign img[10360] = 254;
assign img[10361] = 191;
assign img[10362] = 187;
assign img[10363] = 187;
assign img[10364] = 219;
assign img[10365] = 255;
assign img[10366] = 255;
assign img[10367] = 255;
assign img[10368] = 96;
assign img[10369] = 238;
assign img[10370] = 238;
assign img[10371] = 206;
assign img[10372] = 204;
assign img[10373] = 236;
assign img[10374] = 238;
assign img[10375] = 238;
assign img[10376] = 238;
assign img[10377] = 238;
assign img[10378] = 238;
assign img[10379] = 238;
assign img[10380] = 254;
assign img[10381] = 255;
assign img[10382] = 238;
assign img[10383] = 222;
assign img[10384] = 236;
assign img[10385] = 255;
assign img[10386] = 255;
assign img[10387] = 255;
assign img[10388] = 255;
assign img[10389] = 255;
assign img[10390] = 255;
assign img[10391] = 255;
assign img[10392] = 255;
assign img[10393] = 191;
assign img[10394] = 171;
assign img[10395] = 238;
assign img[10396] = 238;
assign img[10397] = 255;
assign img[10398] = 239;
assign img[10399] = 206;
assign img[10400] = 220;
assign img[10401] = 253;
assign img[10402] = 255;
assign img[10403] = 255;
assign img[10404] = 255;
assign img[10405] = 255;
assign img[10406] = 255;
assign img[10407] = 255;
assign img[10408] = 255;
assign img[10409] = 255;
assign img[10410] = 191;
assign img[10411] = 255;
assign img[10412] = 238;
assign img[10413] = 238;
assign img[10414] = 204;
assign img[10415] = 239;
assign img[10416] = 254;
assign img[10417] = 255;
assign img[10418] = 255;
assign img[10419] = 223;
assign img[10420] = 204;
assign img[10421] = 254;
assign img[10422] = 255;
assign img[10423] = 255;
assign img[10424] = 255;
assign img[10425] = 255;
assign img[10426] = 255;
assign img[10427] = 255;
assign img[10428] = 238;
assign img[10429] = 238;
assign img[10430] = 238;
assign img[10431] = 238;
assign img[10432] = 238;
assign img[10433] = 255;
assign img[10434] = 255;
assign img[10435] = 255;
assign img[10436] = 255;
assign img[10437] = 239;
assign img[10438] = 254;
assign img[10439] = 255;
assign img[10440] = 255;
assign img[10441] = 255;
assign img[10442] = 255;
assign img[10443] = 255;
assign img[10444] = 255;
assign img[10445] = 255;
assign img[10446] = 255;
assign img[10447] = 255;
assign img[10448] = 255;
assign img[10449] = 255;
assign img[10450] = 255;
assign img[10451] = 255;
assign img[10452] = 239;
assign img[10453] = 255;
assign img[10454] = 255;
assign img[10455] = 255;
assign img[10456] = 255;
assign img[10457] = 255;
assign img[10458] = 255;
assign img[10459] = 255;
assign img[10460] = 255;
assign img[10461] = 255;
assign img[10462] = 255;
assign img[10463] = 255;
assign img[10464] = 221;
assign img[10465] = 221;
assign img[10466] = 253;
assign img[10467] = 255;
assign img[10468] = 255;
assign img[10469] = 255;
assign img[10470] = 255;
assign img[10471] = 255;
assign img[10472] = 255;
assign img[10473] = 255;
assign img[10474] = 255;
assign img[10475] = 255;
assign img[10476] = 222;
assign img[10477] = 255;
assign img[10478] = 238;
assign img[10479] = 238;
assign img[10480] = 238;
assign img[10481] = 239;
assign img[10482] = 238;
assign img[10483] = 238;
assign img[10484] = 238;
assign img[10485] = 238;
assign img[10486] = 238;
assign img[10487] = 238;
assign img[10488] = 238;
assign img[10489] = 238;
assign img[10490] = 238;
assign img[10491] = 255;
assign img[10492] = 255;
assign img[10493] = 255;
assign img[10494] = 255;
assign img[10495] = 239;
assign img[10496] = 32;
assign img[10497] = 34;
assign img[10498] = 98;
assign img[10499] = 247;
assign img[10500] = 255;
assign img[10501] = 255;
assign img[10502] = 255;
assign img[10503] = 223;
assign img[10504] = 253;
assign img[10505] = 255;
assign img[10506] = 255;
assign img[10507] = 239;
assign img[10508] = 206;
assign img[10509] = 238;
assign img[10510] = 174;
assign img[10511] = 138;
assign img[10512] = 200;
assign img[10513] = 205;
assign img[10514] = 236;
assign img[10515] = 255;
assign img[10516] = 221;
assign img[10517] = 221;
assign img[10518] = 221;
assign img[10519] = 253;
assign img[10520] = 255;
assign img[10521] = 255;
assign img[10522] = 239;
assign img[10523] = 238;
assign img[10524] = 238;
assign img[10525] = 255;
assign img[10526] = 255;
assign img[10527] = 191;
assign img[10528] = 187;
assign img[10529] = 251;
assign img[10530] = 255;
assign img[10531] = 255;
assign img[10532] = 223;
assign img[10533] = 255;
assign img[10534] = 255;
assign img[10535] = 255;
assign img[10536] = 238;
assign img[10537] = 238;
assign img[10538] = 238;
assign img[10539] = 255;
assign img[10540] = 238;
assign img[10541] = 239;
assign img[10542] = 238;
assign img[10543] = 238;
assign img[10544] = 238;
assign img[10545] = 238;
assign img[10546] = 238;
assign img[10547] = 238;
assign img[10548] = 254;
assign img[10549] = 239;
assign img[10550] = 238;
assign img[10551] = 238;
assign img[10552] = 238;
assign img[10553] = 255;
assign img[10554] = 255;
assign img[10555] = 255;
assign img[10556] = 238;
assign img[10557] = 255;
assign img[10558] = 238;
assign img[10559] = 255;
assign img[10560] = 255;
assign img[10561] = 255;
assign img[10562] = 239;
assign img[10563] = 238;
assign img[10564] = 238;
assign img[10565] = 238;
assign img[10566] = 238;
assign img[10567] = 238;
assign img[10568] = 238;
assign img[10569] = 238;
assign img[10570] = 238;
assign img[10571] = 238;
assign img[10572] = 238;
assign img[10573] = 238;
assign img[10574] = 238;
assign img[10575] = 238;
assign img[10576] = 238;
assign img[10577] = 254;
assign img[10578] = 238;
assign img[10579] = 238;
assign img[10580] = 238;
assign img[10581] = 254;
assign img[10582] = 255;
assign img[10583] = 255;
assign img[10584] = 239;
assign img[10585] = 238;
assign img[10586] = 238;
assign img[10587] = 206;
assign img[10588] = 254;
assign img[10589] = 255;
assign img[10590] = 255;
assign img[10591] = 191;
assign img[10592] = 255;
assign img[10593] = 255;
assign img[10594] = 255;
assign img[10595] = 255;
assign img[10596] = 255;
assign img[10597] = 255;
assign img[10598] = 206;
assign img[10599] = 204;
assign img[10600] = 236;
assign img[10601] = 255;
assign img[10602] = 204;
assign img[10603] = 221;
assign img[10604] = 204;
assign img[10605] = 253;
assign img[10606] = 238;
assign img[10607] = 238;
assign img[10608] = 220;
assign img[10609] = 157;
assign img[10610] = 249;
assign img[10611] = 255;
assign img[10612] = 255;
assign img[10613] = 255;
assign img[10614] = 255;
assign img[10615] = 255;
assign img[10616] = 223;
assign img[10617] = 255;
assign img[10618] = 187;
assign img[10619] = 251;
assign img[10620] = 255;
assign img[10621] = 255;
assign img[10622] = 255;
assign img[10623] = 255;
assign img[10624] = 32;
assign img[10625] = 255;
assign img[10626] = 255;
assign img[10627] = 255;
assign img[10628] = 253;
assign img[10629] = 204;
assign img[10630] = 204;
assign img[10631] = 238;
assign img[10632] = 238;
assign img[10633] = 255;
assign img[10634] = 255;
assign img[10635] = 255;
assign img[10636] = 205;
assign img[10637] = 238;
assign img[10638] = 238;
assign img[10639] = 239;
assign img[10640] = 238;
assign img[10641] = 238;
assign img[10642] = 254;
assign img[10643] = 255;
assign img[10644] = 187;
assign img[10645] = 255;
assign img[10646] = 254;
assign img[10647] = 255;
assign img[10648] = 254;
assign img[10649] = 238;
assign img[10650] = 254;
assign img[10651] = 255;
assign img[10652] = 255;
assign img[10653] = 255;
assign img[10654] = 255;
assign img[10655] = 255;
assign img[10656] = 255;
assign img[10657] = 255;
assign img[10658] = 255;
assign img[10659] = 255;
assign img[10660] = 255;
assign img[10661] = 255;
assign img[10662] = 255;
assign img[10663] = 255;
assign img[10664] = 254;
assign img[10665] = 255;
assign img[10666] = 223;
assign img[10667] = 204;
assign img[10668] = 236;
assign img[10669] = 238;
assign img[10670] = 238;
assign img[10671] = 255;
assign img[10672] = 255;
assign img[10673] = 255;
assign img[10674] = 255;
assign img[10675] = 255;
assign img[10676] = 255;
assign img[10677] = 255;
assign img[10678] = 255;
assign img[10679] = 255;
assign img[10680] = 191;
assign img[10681] = 187;
assign img[10682] = 219;
assign img[10683] = 255;
assign img[10684] = 255;
assign img[10685] = 239;
assign img[10686] = 238;
assign img[10687] = 255;
assign img[10688] = 255;
assign img[10689] = 255;
assign img[10690] = 255;
assign img[10691] = 255;
assign img[10692] = 255;
assign img[10693] = 255;
assign img[10694] = 205;
assign img[10695] = 238;
assign img[10696] = 238;
assign img[10697] = 255;
assign img[10698] = 255;
assign img[10699] = 255;
assign img[10700] = 255;
assign img[10701] = 255;
assign img[10702] = 255;
assign img[10703] = 255;
assign img[10704] = 255;
assign img[10705] = 255;
assign img[10706] = 255;
assign img[10707] = 255;
assign img[10708] = 223;
assign img[10709] = 204;
assign img[10710] = 236;
assign img[10711] = 238;
assign img[10712] = 254;
assign img[10713] = 255;
assign img[10714] = 255;
assign img[10715] = 255;
assign img[10716] = 255;
assign img[10717] = 255;
assign img[10718] = 255;
assign img[10719] = 255;
assign img[10720] = 187;
assign img[10721] = 139;
assign img[10722] = 248;
assign img[10723] = 255;
assign img[10724] = 255;
assign img[10725] = 255;
assign img[10726] = 255;
assign img[10727] = 255;
assign img[10728] = 255;
assign img[10729] = 255;
assign img[10730] = 255;
assign img[10731] = 255;
assign img[10732] = 255;
assign img[10733] = 255;
assign img[10734] = 255;
assign img[10735] = 255;
assign img[10736] = 239;
assign img[10737] = 238;
assign img[10738] = 238;
assign img[10739] = 239;
assign img[10740] = 238;
assign img[10741] = 238;
assign img[10742] = 238;
assign img[10743] = 238;
assign img[10744] = 238;
assign img[10745] = 255;
assign img[10746] = 239;
assign img[10747] = 223;
assign img[10748] = 221;
assign img[10749] = 253;
assign img[10750] = 223;
assign img[10751] = 221;
assign img[10752] = 96;
assign img[10753] = 255;
assign img[10754] = 255;
assign img[10755] = 223;
assign img[10756] = 221;
assign img[10757] = 221;
assign img[10758] = 221;
assign img[10759] = 239;
assign img[10760] = 238;
assign img[10761] = 238;
assign img[10762] = 254;
assign img[10763] = 255;
assign img[10764] = 155;
assign img[10765] = 153;
assign img[10766] = 221;
assign img[10767] = 221;
assign img[10768] = 221;
assign img[10769] = 207;
assign img[10770] = 238;
assign img[10771] = 238;
assign img[10772] = 186;
assign img[10773] = 255;
assign img[10774] = 255;
assign img[10775] = 255;
assign img[10776] = 255;
assign img[10777] = 239;
assign img[10778] = 238;
assign img[10779] = 238;
assign img[10780] = 238;
assign img[10781] = 254;
assign img[10782] = 238;
assign img[10783] = 206;
assign img[10784] = 204;
assign img[10785] = 255;
assign img[10786] = 239;
assign img[10787] = 254;
assign img[10788] = 255;
assign img[10789] = 255;
assign img[10790] = 238;
assign img[10791] = 238;
assign img[10792] = 238;
assign img[10793] = 255;
assign img[10794] = 255;
assign img[10795] = 255;
assign img[10796] = 255;
assign img[10797] = 255;
assign img[10798] = 238;
assign img[10799] = 255;
assign img[10800] = 255;
assign img[10801] = 255;
assign img[10802] = 255;
assign img[10803] = 255;
assign img[10804] = 255;
assign img[10805] = 255;
assign img[10806] = 238;
assign img[10807] = 238;
assign img[10808] = 238;
assign img[10809] = 238;
assign img[10810] = 206;
assign img[10811] = 204;
assign img[10812] = 236;
assign img[10813] = 238;
assign img[10814] = 238;
assign img[10815] = 255;
assign img[10816] = 255;
assign img[10817] = 255;
assign img[10818] = 255;
assign img[10819] = 255;
assign img[10820] = 255;
assign img[10821] = 255;
assign img[10822] = 238;
assign img[10823] = 238;
assign img[10824] = 255;
assign img[10825] = 254;
assign img[10826] = 238;
assign img[10827] = 238;
assign img[10828] = 238;
assign img[10829] = 238;
assign img[10830] = 238;
assign img[10831] = 238;
assign img[10832] = 238;
assign img[10833] = 254;
assign img[10834] = 255;
assign img[10835] = 254;
assign img[10836] = 255;
assign img[10837] = 255;
assign img[10838] = 255;
assign img[10839] = 255;
assign img[10840] = 255;
assign img[10841] = 255;
assign img[10842] = 239;
assign img[10843] = 238;
assign img[10844] = 254;
assign img[10845] = 255;
assign img[10846] = 255;
assign img[10847] = 239;
assign img[10848] = 238;
assign img[10849] = 238;
assign img[10850] = 238;
assign img[10851] = 238;
assign img[10852] = 238;
assign img[10853] = 238;
assign img[10854] = 206;
assign img[10855] = 238;
assign img[10856] = 238;
assign img[10857] = 238;
assign img[10858] = 238;
assign img[10859] = 206;
assign img[10860] = 254;
assign img[10861] = 255;
assign img[10862] = 223;
assign img[10863] = 221;
assign img[10864] = 255;
assign img[10865] = 255;
assign img[10866] = 221;
assign img[10867] = 221;
assign img[10868] = 253;
assign img[10869] = 255;
assign img[10870] = 255;
assign img[10871] = 255;
assign img[10872] = 255;
assign img[10873] = 239;
assign img[10874] = 206;
assign img[10875] = 206;
assign img[10876] = 204;
assign img[10877] = 252;
assign img[10878] = 239;
assign img[10879] = 238;
assign img[10880] = 96;
assign img[10881] = 239;
assign img[10882] = 238;
assign img[10883] = 255;
assign img[10884] = 239;
assign img[10885] = 238;
assign img[10886] = 238;
assign img[10887] = 254;
assign img[10888] = 239;
assign img[10889] = 238;
assign img[10890] = 238;
assign img[10891] = 238;
assign img[10892] = 254;
assign img[10893] = 255;
assign img[10894] = 223;
assign img[10895] = 221;
assign img[10896] = 221;
assign img[10897] = 255;
assign img[10898] = 255;
assign img[10899] = 239;
assign img[10900] = 238;
assign img[10901] = 238;
assign img[10902] = 238;
assign img[10903] = 255;
assign img[10904] = 255;
assign img[10905] = 239;
assign img[10906] = 238;
assign img[10907] = 238;
assign img[10908] = 238;
assign img[10909] = 255;
assign img[10910] = 239;
assign img[10911] = 206;
assign img[10912] = 254;
assign img[10913] = 255;
assign img[10914] = 255;
assign img[10915] = 255;
assign img[10916] = 239;
assign img[10917] = 255;
assign img[10918] = 255;
assign img[10919] = 255;
assign img[10920] = 255;
assign img[10921] = 255;
assign img[10922] = 255;
assign img[10923] = 255;
assign img[10924] = 255;
assign img[10925] = 238;
assign img[10926] = 238;
assign img[10927] = 255;
assign img[10928] = 255;
assign img[10929] = 255;
assign img[10930] = 255;
assign img[10931] = 255;
assign img[10932] = 255;
assign img[10933] = 255;
assign img[10934] = 255;
assign img[10935] = 255;
assign img[10936] = 255;
assign img[10937] = 223;
assign img[10938] = 238;
assign img[10939] = 238;
assign img[10940] = 238;
assign img[10941] = 238;
assign img[10942] = 238;
assign img[10943] = 255;
assign img[10944] = 255;
assign img[10945] = 255;
assign img[10946] = 255;
assign img[10947] = 255;
assign img[10948] = 255;
assign img[10949] = 255;
assign img[10950] = 139;
assign img[10951] = 238;
assign img[10952] = 238;
assign img[10953] = 238;
assign img[10954] = 254;
assign img[10955] = 239;
assign img[10956] = 238;
assign img[10957] = 238;
assign img[10958] = 238;
assign img[10959] = 255;
assign img[10960] = 223;
assign img[10961] = 255;
assign img[10962] = 255;
assign img[10963] = 239;
assign img[10964] = 186;
assign img[10965] = 239;
assign img[10966] = 238;
assign img[10967] = 238;
assign img[10968] = 206;
assign img[10969] = 255;
assign img[10970] = 255;
assign img[10971] = 255;
assign img[10972] = 255;
assign img[10973] = 255;
assign img[10974] = 255;
assign img[10975] = 191;
assign img[10976] = 187;
assign img[10977] = 187;
assign img[10978] = 251;
assign img[10979] = 255;
assign img[10980] = 255;
assign img[10981] = 239;
assign img[10982] = 206;
assign img[10983] = 254;
assign img[10984] = 238;
assign img[10985] = 238;
assign img[10986] = 238;
assign img[10987] = 238;
assign img[10988] = 206;
assign img[10989] = 204;
assign img[10990] = 204;
assign img[10991] = 255;
assign img[10992] = 223;
assign img[10993] = 221;
assign img[10994] = 253;
assign img[10995] = 255;
assign img[10996] = 223;
assign img[10997] = 221;
assign img[10998] = 221;
assign img[10999] = 255;
assign img[11000] = 254;
assign img[11001] = 255;
assign img[11002] = 255;
assign img[11003] = 255;
assign img[11004] = 238;
assign img[11005] = 238;
assign img[11006] = 206;
assign img[11007] = 238;
assign img[11008] = 0;
assign img[11009] = 196;
assign img[11010] = 252;
assign img[11011] = 223;
assign img[11012] = 221;
assign img[11013] = 221;
assign img[11014] = 137;
assign img[11015] = 234;
assign img[11016] = 238;
assign img[11017] = 238;
assign img[11018] = 254;
assign img[11019] = 223;
assign img[11020] = 221;
assign img[11021] = 253;
assign img[11022] = 255;
assign img[11023] = 239;
assign img[11024] = 238;
assign img[11025] = 222;
assign img[11026] = 221;
assign img[11027] = 223;
assign img[11028] = 236;
assign img[11029] = 255;
assign img[11030] = 255;
assign img[11031] = 255;
assign img[11032] = 255;
assign img[11033] = 239;
assign img[11034] = 254;
assign img[11035] = 255;
assign img[11036] = 255;
assign img[11037] = 255;
assign img[11038] = 255;
assign img[11039] = 191;
assign img[11040] = 187;
assign img[11041] = 251;
assign img[11042] = 255;
assign img[11043] = 255;
assign img[11044] = 255;
assign img[11045] = 255;
assign img[11046] = 255;
assign img[11047] = 255;
assign img[11048] = 255;
assign img[11049] = 255;
assign img[11050] = 255;
assign img[11051] = 255;
assign img[11052] = 255;
assign img[11053] = 255;
assign img[11054] = 254;
assign img[11055] = 255;
assign img[11056] = 255;
assign img[11057] = 255;
assign img[11058] = 255;
assign img[11059] = 255;
assign img[11060] = 191;
assign img[11061] = 255;
assign img[11062] = 255;
assign img[11063] = 255;
assign img[11064] = 255;
assign img[11065] = 255;
assign img[11066] = 239;
assign img[11067] = 238;
assign img[11068] = 238;
assign img[11069] = 255;
assign img[11070] = 239;
assign img[11071] = 255;
assign img[11072] = 255;
assign img[11073] = 255;
assign img[11074] = 255;
assign img[11075] = 255;
assign img[11076] = 255;
assign img[11077] = 239;
assign img[11078] = 254;
assign img[11079] = 255;
assign img[11080] = 255;
assign img[11081] = 255;
assign img[11082] = 255;
assign img[11083] = 255;
assign img[11084] = 255;
assign img[11085] = 255;
assign img[11086] = 255;
assign img[11087] = 255;
assign img[11088] = 255;
assign img[11089] = 255;
assign img[11090] = 255;
assign img[11091] = 255;
assign img[11092] = 223;
assign img[11093] = 255;
assign img[11094] = 255;
assign img[11095] = 255;
assign img[11096] = 255;
assign img[11097] = 255;
assign img[11098] = 223;
assign img[11099] = 255;
assign img[11100] = 255;
assign img[11101] = 255;
assign img[11102] = 255;
assign img[11103] = 191;
assign img[11104] = 255;
assign img[11105] = 239;
assign img[11106] = 254;
assign img[11107] = 255;
assign img[11108] = 255;
assign img[11109] = 255;
assign img[11110] = 255;
assign img[11111] = 255;
assign img[11112] = 254;
assign img[11113] = 238;
assign img[11114] = 204;
assign img[11115] = 238;
assign img[11116] = 206;
assign img[11117] = 238;
assign img[11118] = 206;
assign img[11119] = 255;
assign img[11120] = 255;
assign img[11121] = 238;
assign img[11122] = 254;
assign img[11123] = 255;
assign img[11124] = 221;
assign img[11125] = 221;
assign img[11126] = 253;
assign img[11127] = 255;
assign img[11128] = 255;
assign img[11129] = 255;
assign img[11130] = 238;
assign img[11131] = 238;
assign img[11132] = 222;
assign img[11133] = 255;
assign img[11134] = 255;
assign img[11135] = 239;
assign img[11136] = 96;
assign img[11137] = 206;
assign img[11138] = 252;
assign img[11139] = 239;
assign img[11140] = 238;
assign img[11141] = 238;
assign img[11142] = 206;
assign img[11143] = 238;
assign img[11144] = 238;
assign img[11145] = 238;
assign img[11146] = 238;
assign img[11147] = 255;
assign img[11148] = 157;
assign img[11149] = 187;
assign img[11150] = 251;
assign img[11151] = 255;
assign img[11152] = 239;
assign img[11153] = 238;
assign img[11154] = 238;
assign img[11155] = 238;
assign img[11156] = 220;
assign img[11157] = 255;
assign img[11158] = 255;
assign img[11159] = 255;
assign img[11160] = 238;
assign img[11161] = 255;
assign img[11162] = 255;
assign img[11163] = 255;
assign img[11164] = 255;
assign img[11165] = 255;
assign img[11166] = 255;
assign img[11167] = 223;
assign img[11168] = 204;
assign img[11169] = 236;
assign img[11170] = 238;
assign img[11171] = 255;
assign img[11172] = 223;
assign img[11173] = 255;
assign img[11174] = 238;
assign img[11175] = 255;
assign img[11176] = 238;
assign img[11177] = 238;
assign img[11178] = 238;
assign img[11179] = 238;
assign img[11180] = 238;
assign img[11181] = 238;
assign img[11182] = 238;
assign img[11183] = 206;
assign img[11184] = 238;
assign img[11185] = 206;
assign img[11186] = 236;
assign img[11187] = 238;
assign img[11188] = 206;
assign img[11189] = 255;
assign img[11190] = 255;
assign img[11191] = 255;
assign img[11192] = 255;
assign img[11193] = 255;
assign img[11194] = 255;
assign img[11195] = 255;
assign img[11196] = 238;
assign img[11197] = 255;
assign img[11198] = 254;
assign img[11199] = 255;
assign img[11200] = 254;
assign img[11201] = 255;
assign img[11202] = 238;
assign img[11203] = 255;
assign img[11204] = 254;
assign img[11205] = 255;
assign img[11206] = 238;
assign img[11207] = 238;
assign img[11208] = 238;
assign img[11209] = 238;
assign img[11210] = 254;
assign img[11211] = 223;
assign img[11212] = 255;
assign img[11213] = 255;
assign img[11214] = 255;
assign img[11215] = 255;
assign img[11216] = 255;
assign img[11217] = 255;
assign img[11218] = 239;
assign img[11219] = 239;
assign img[11220] = 239;
assign img[11221] = 238;
assign img[11222] = 238;
assign img[11223] = 238;
assign img[11224] = 238;
assign img[11225] = 238;
assign img[11226] = 238;
assign img[11227] = 206;
assign img[11228] = 252;
assign img[11229] = 255;
assign img[11230] = 255;
assign img[11231] = 223;
assign img[11232] = 221;
assign img[11233] = 205;
assign img[11234] = 236;
assign img[11235] = 238;
assign img[11236] = 238;
assign img[11237] = 206;
assign img[11238] = 236;
assign img[11239] = 254;
assign img[11240] = 238;
assign img[11241] = 254;
assign img[11242] = 238;
assign img[11243] = 255;
assign img[11244] = 223;
assign img[11245] = 255;
assign img[11246] = 255;
assign img[11247] = 239;
assign img[11248] = 254;
assign img[11249] = 255;
assign img[11250] = 255;
assign img[11251] = 191;
assign img[11252] = 155;
assign img[11253] = 255;
assign img[11254] = 223;
assign img[11255] = 253;
assign img[11256] = 255;
assign img[11257] = 255;
assign img[11258] = 255;
assign img[11259] = 255;
assign img[11260] = 221;
assign img[11261] = 255;
assign img[11262] = 223;
assign img[11263] = 255;
assign img[11264] = 96;
assign img[11265] = 223;
assign img[11266] = 253;
assign img[11267] = 255;
assign img[11268] = 223;
assign img[11269] = 253;
assign img[11270] = 223;
assign img[11271] = 253;
assign img[11272] = 255;
assign img[11273] = 255;
assign img[11274] = 255;
assign img[11275] = 255;
assign img[11276] = 255;
assign img[11277] = 255;
assign img[11278] = 191;
assign img[11279] = 187;
assign img[11280] = 217;
assign img[11281] = 253;
assign img[11282] = 255;
assign img[11283] = 255;
assign img[11284] = 221;
assign img[11285] = 255;
assign img[11286] = 223;
assign img[11287] = 255;
assign img[11288] = 255;
assign img[11289] = 255;
assign img[11290] = 205;
assign img[11291] = 238;
assign img[11292] = 238;
assign img[11293] = 255;
assign img[11294] = 223;
assign img[11295] = 191;
assign img[11296] = 155;
assign img[11297] = 255;
assign img[11298] = 255;
assign img[11299] = 255;
assign img[11300] = 255;
assign img[11301] = 255;
assign img[11302] = 255;
assign img[11303] = 255;
assign img[11304] = 255;
assign img[11305] = 255;
assign img[11306] = 255;
assign img[11307] = 239;
assign img[11308] = 238;
assign img[11309] = 238;
assign img[11310] = 238;
assign img[11311] = 238;
assign img[11312] = 254;
assign img[11313] = 255;
assign img[11314] = 239;
assign img[11315] = 254;
assign img[11316] = 255;
assign img[11317] = 255;
assign img[11318] = 255;
assign img[11319] = 255;
assign img[11320] = 255;
assign img[11321] = 255;
assign img[11322] = 223;
assign img[11323] = 255;
assign img[11324] = 255;
assign img[11325] = 255;
assign img[11326] = 238;
assign img[11327] = 255;
assign img[11328] = 255;
assign img[11329] = 255;
assign img[11330] = 239;
assign img[11331] = 238;
assign img[11332] = 238;
assign img[11333] = 206;
assign img[11334] = 238;
assign img[11335] = 238;
assign img[11336] = 238;
assign img[11337] = 255;
assign img[11338] = 255;
assign img[11339] = 223;
assign img[11340] = 255;
assign img[11341] = 255;
assign img[11342] = 238;
assign img[11343] = 255;
assign img[11344] = 239;
assign img[11345] = 238;
assign img[11346] = 238;
assign img[11347] = 255;
assign img[11348] = 239;
assign img[11349] = 254;
assign img[11350] = 238;
assign img[11351] = 255;
assign img[11352] = 255;
assign img[11353] = 255;
assign img[11354] = 255;
assign img[11355] = 239;
assign img[11356] = 254;
assign img[11357] = 255;
assign img[11358] = 255;
assign img[11359] = 223;
assign img[11360] = 189;
assign img[11361] = 155;
assign img[11362] = 249;
assign img[11363] = 255;
assign img[11364] = 255;
assign img[11365] = 255;
assign img[11366] = 206;
assign img[11367] = 238;
assign img[11368] = 255;
assign img[11369] = 255;
assign img[11370] = 255;
assign img[11371] = 255;
assign img[11372] = 255;
assign img[11373] = 255;
assign img[11374] = 255;
assign img[11375] = 239;
assign img[11376] = 238;
assign img[11377] = 174;
assign img[11378] = 170;
assign img[11379] = 255;
assign img[11380] = 255;
assign img[11381] = 239;
assign img[11382] = 238;
assign img[11383] = 238;
assign img[11384] = 238;
assign img[11385] = 238;
assign img[11386] = 204;
assign img[11387] = 204;
assign img[11388] = 236;
assign img[11389] = 238;
assign img[11390] = 238;
assign img[11391] = 238;
assign img[11392] = 64;
assign img[11393] = 68;
assign img[11394] = 116;
assign img[11395] = 255;
assign img[11396] = 255;
assign img[11397] = 223;
assign img[11398] = 221;
assign img[11399] = 255;
assign img[11400] = 255;
assign img[11401] = 255;
assign img[11402] = 255;
assign img[11403] = 255;
assign img[11404] = 255;
assign img[11405] = 255;
assign img[11406] = 223;
assign img[11407] = 221;
assign img[11408] = 236;
assign img[11409] = 238;
assign img[11410] = 254;
assign img[11411] = 223;
assign img[11412] = 236;
assign img[11413] = 254;
assign img[11414] = 204;
assign img[11415] = 238;
assign img[11416] = 238;
assign img[11417] = 207;
assign img[11418] = 204;
assign img[11419] = 204;
assign img[11420] = 236;
assign img[11421] = 255;
assign img[11422] = 223;
assign img[11423] = 221;
assign img[11424] = 221;
assign img[11425] = 253;
assign img[11426] = 255;
assign img[11427] = 255;
assign img[11428] = 255;
assign img[11429] = 255;
assign img[11430] = 255;
assign img[11431] = 207;
assign img[11432] = 236;
assign img[11433] = 238;
assign img[11434] = 254;
assign img[11435] = 255;
assign img[11436] = 239;
assign img[11437] = 238;
assign img[11438] = 238;
assign img[11439] = 238;
assign img[11440] = 254;
assign img[11441] = 255;
assign img[11442] = 239;
assign img[11443] = 238;
assign img[11444] = 238;
assign img[11445] = 254;
assign img[11446] = 239;
assign img[11447] = 239;
assign img[11448] = 238;
assign img[11449] = 239;
assign img[11450] = 254;
assign img[11451] = 255;
assign img[11452] = 255;
assign img[11453] = 223;
assign img[11454] = 221;
assign img[11455] = 255;
assign img[11456] = 255;
assign img[11457] = 255;
assign img[11458] = 238;
assign img[11459] = 238;
assign img[11460] = 255;
assign img[11461] = 223;
assign img[11462] = 253;
assign img[11463] = 255;
assign img[11464] = 255;
assign img[11465] = 255;
assign img[11466] = 255;
assign img[11467] = 255;
assign img[11468] = 255;
assign img[11469] = 255;
assign img[11470] = 255;
assign img[11471] = 255;
assign img[11472] = 255;
assign img[11473] = 255;
assign img[11474] = 255;
assign img[11475] = 255;
assign img[11476] = 255;
assign img[11477] = 255;
assign img[11478] = 255;
assign img[11479] = 255;
assign img[11480] = 239;
assign img[11481] = 238;
assign img[11482] = 206;
assign img[11483] = 238;
assign img[11484] = 254;
assign img[11485] = 255;
assign img[11486] = 255;
assign img[11487] = 239;
assign img[11488] = 204;
assign img[11489] = 204;
assign img[11490] = 252;
assign img[11491] = 255;
assign img[11492] = 255;
assign img[11493] = 255;
assign img[11494] = 239;
assign img[11495] = 238;
assign img[11496] = 238;
assign img[11497] = 239;
assign img[11498] = 238;
assign img[11499] = 238;
assign img[11500] = 238;
assign img[11501] = 254;
assign img[11502] = 255;
assign img[11503] = 255;
assign img[11504] = 206;
assign img[11505] = 220;
assign img[11506] = 236;
assign img[11507] = 255;
assign img[11508] = 204;
assign img[11509] = 255;
assign img[11510] = 254;
assign img[11511] = 255;
assign img[11512] = 254;
assign img[11513] = 238;
assign img[11514] = 220;
assign img[11515] = 237;
assign img[11516] = 238;
assign img[11517] = 254;
assign img[11518] = 255;
assign img[11519] = 223;
assign img[11520] = 96;
assign img[11521] = 223;
assign img[11522] = 205;
assign img[11523] = 220;
assign img[11524] = 169;
assign img[11525] = 138;
assign img[11526] = 184;
assign img[11527] = 239;
assign img[11528] = 238;
assign img[11529] = 238;
assign img[11530] = 238;
assign img[11531] = 238;
assign img[11532] = 238;
assign img[11533] = 238;
assign img[11534] = 170;
assign img[11535] = 170;
assign img[11536] = 238;
assign img[11537] = 255;
assign img[11538] = 255;
assign img[11539] = 239;
assign img[11540] = 238;
assign img[11541] = 204;
assign img[11542] = 204;
assign img[11543] = 236;
assign img[11544] = 238;
assign img[11545] = 207;
assign img[11546] = 204;
assign img[11547] = 238;
assign img[11548] = 238;
assign img[11549] = 254;
assign img[11550] = 255;
assign img[11551] = 238;
assign img[11552] = 254;
assign img[11553] = 255;
assign img[11554] = 255;
assign img[11555] = 255;
assign img[11556] = 239;
assign img[11557] = 238;
assign img[11558] = 238;
assign img[11559] = 239;
assign img[11560] = 238;
assign img[11561] = 238;
assign img[11562] = 254;
assign img[11563] = 255;
assign img[11564] = 255;
assign img[11565] = 239;
assign img[11566] = 238;
assign img[11567] = 238;
assign img[11568] = 238;
assign img[11569] = 238;
assign img[11570] = 238;
assign img[11571] = 255;
assign img[11572] = 255;
assign img[11573] = 255;
assign img[11574] = 255;
assign img[11575] = 255;
assign img[11576] = 255;
assign img[11577] = 255;
assign img[11578] = 255;
assign img[11579] = 239;
assign img[11580] = 238;
assign img[11581] = 238;
assign img[11582] = 254;
assign img[11583] = 255;
assign img[11584] = 255;
assign img[11585] = 255;
assign img[11586] = 255;
assign img[11587] = 255;
assign img[11588] = 255;
assign img[11589] = 255;
assign img[11590] = 255;
assign img[11591] = 255;
assign img[11592] = 255;
assign img[11593] = 255;
assign img[11594] = 255;
assign img[11595] = 255;
assign img[11596] = 191;
assign img[11597] = 255;
assign img[11598] = 254;
assign img[11599] = 255;
assign img[11600] = 223;
assign img[11601] = 255;
assign img[11602] = 239;
assign img[11603] = 238;
assign img[11604] = 238;
assign img[11605] = 238;
assign img[11606] = 238;
assign img[11607] = 238;
assign img[11608] = 238;
assign img[11609] = 238;
assign img[11610] = 238;
assign img[11611] = 238;
assign img[11612] = 254;
assign img[11613] = 255;
assign img[11614] = 255;
assign img[11615] = 207;
assign img[11616] = 204;
assign img[11617] = 238;
assign img[11618] = 238;
assign img[11619] = 238;
assign img[11620] = 238;
assign img[11621] = 255;
assign img[11622] = 207;
assign img[11623] = 220;
assign img[11624] = 253;
assign img[11625] = 223;
assign img[11626] = 253;
assign img[11627] = 255;
assign img[11628] = 238;
assign img[11629] = 238;
assign img[11630] = 238;
assign img[11631] = 255;
assign img[11632] = 255;
assign img[11633] = 255;
assign img[11634] = 238;
assign img[11635] = 238;
assign img[11636] = 254;
assign img[11637] = 255;
assign img[11638] = 238;
assign img[11639] = 238;
assign img[11640] = 238;
assign img[11641] = 206;
assign img[11642] = 204;
assign img[11643] = 204;
assign img[11644] = 204;
assign img[11645] = 239;
assign img[11646] = 238;
assign img[11647] = 238;
assign img[11648] = 96;
assign img[11649] = 223;
assign img[11650] = 253;
assign img[11651] = 239;
assign img[11652] = 170;
assign img[11653] = 255;
assign img[11654] = 255;
assign img[11655] = 255;
assign img[11656] = 255;
assign img[11657] = 255;
assign img[11658] = 255;
assign img[11659] = 255;
assign img[11660] = 157;
assign img[11661] = 253;
assign img[11662] = 191;
assign img[11663] = 223;
assign img[11664] = 221;
assign img[11665] = 253;
assign img[11666] = 255;
assign img[11667] = 239;
assign img[11668] = 254;
assign img[11669] = 255;
assign img[11670] = 239;
assign img[11671] = 255;
assign img[11672] = 255;
assign img[11673] = 239;
assign img[11674] = 238;
assign img[11675] = 238;
assign img[11676] = 238;
assign img[11677] = 255;
assign img[11678] = 255;
assign img[11679] = 239;
assign img[11680] = 238;
assign img[11681] = 238;
assign img[11682] = 238;
assign img[11683] = 255;
assign img[11684] = 255;
assign img[11685] = 255;
assign img[11686] = 255;
assign img[11687] = 239;
assign img[11688] = 238;
assign img[11689] = 238;
assign img[11690] = 254;
assign img[11691] = 255;
assign img[11692] = 255;
assign img[11693] = 255;
assign img[11694] = 255;
assign img[11695] = 223;
assign img[11696] = 255;
assign img[11697] = 255;
assign img[11698] = 255;
assign img[11699] = 255;
assign img[11700] = 255;
assign img[11701] = 255;
assign img[11702] = 255;
assign img[11703] = 255;
assign img[11704] = 255;
assign img[11705] = 255;
assign img[11706] = 255;
assign img[11707] = 255;
assign img[11708] = 255;
assign img[11709] = 207;
assign img[11710] = 238;
assign img[11711] = 255;
assign img[11712] = 255;
assign img[11713] = 255;
assign img[11714] = 223;
assign img[11715] = 255;
assign img[11716] = 255;
assign img[11717] = 223;
assign img[11718] = 205;
assign img[11719] = 238;
assign img[11720] = 238;
assign img[11721] = 238;
assign img[11722] = 238;
assign img[11723] = 238;
assign img[11724] = 238;
assign img[11725] = 255;
assign img[11726] = 238;
assign img[11727] = 255;
assign img[11728] = 255;
assign img[11729] = 255;
assign img[11730] = 255;
assign img[11731] = 255;
assign img[11732] = 255;
assign img[11733] = 255;
assign img[11734] = 255;
assign img[11735] = 255;
assign img[11736] = 223;
assign img[11737] = 221;
assign img[11738] = 253;
assign img[11739] = 255;
assign img[11740] = 255;
assign img[11741] = 255;
assign img[11742] = 255;
assign img[11743] = 255;
assign img[11744] = 221;
assign img[11745] = 221;
assign img[11746] = 253;
assign img[11747] = 255;
assign img[11748] = 255;
assign img[11749] = 207;
assign img[11750] = 204;
assign img[11751] = 253;
assign img[11752] = 255;
assign img[11753] = 255;
assign img[11754] = 238;
assign img[11755] = 238;
assign img[11756] = 255;
assign img[11757] = 255;
assign img[11758] = 254;
assign img[11759] = 239;
assign img[11760] = 255;
assign img[11761] = 157;
assign img[11762] = 249;
assign img[11763] = 159;
assign img[11764] = 137;
assign img[11765] = 238;
assign img[11766] = 238;
assign img[11767] = 238;
assign img[11768] = 238;
assign img[11769] = 255;
assign img[11770] = 255;
assign img[11771] = 255;
assign img[11772] = 255;
assign img[11773] = 255;
assign img[11774] = 255;
assign img[11775] = 255;
assign img[11776] = 96;
assign img[11777] = 206;
assign img[11778] = 252;
assign img[11779] = 223;
assign img[11780] = 205;
assign img[11781] = 204;
assign img[11782] = 220;
assign img[11783] = 253;
assign img[11784] = 254;
assign img[11785] = 255;
assign img[11786] = 206;
assign img[11787] = 204;
assign img[11788] = 204;
assign img[11789] = 204;
assign img[11790] = 204;
assign img[11791] = 204;
assign img[11792] = 236;
assign img[11793] = 238;
assign img[11794] = 254;
assign img[11795] = 205;
assign img[11796] = 236;
assign img[11797] = 238;
assign img[11798] = 222;
assign img[11799] = 255;
assign img[11800] = 255;
assign img[11801] = 255;
assign img[11802] = 238;
assign img[11803] = 238;
assign img[11804] = 238;
assign img[11805] = 238;
assign img[11806] = 238;
assign img[11807] = 174;
assign img[11808] = 238;
assign img[11809] = 238;
assign img[11810] = 238;
assign img[11811] = 238;
assign img[11812] = 238;
assign img[11813] = 238;
assign img[11814] = 254;
assign img[11815] = 255;
assign img[11816] = 255;
assign img[11817] = 255;
assign img[11818] = 255;
assign img[11819] = 255;
assign img[11820] = 238;
assign img[11821] = 254;
assign img[11822] = 255;
assign img[11823] = 255;
assign img[11824] = 238;
assign img[11825] = 238;
assign img[11826] = 238;
assign img[11827] = 238;
assign img[11828] = 238;
assign img[11829] = 254;
assign img[11830] = 238;
assign img[11831] = 255;
assign img[11832] = 238;
assign img[11833] = 255;
assign img[11834] = 206;
assign img[11835] = 238;
assign img[11836] = 254;
assign img[11837] = 223;
assign img[11838] = 221;
assign img[11839] = 255;
assign img[11840] = 255;
assign img[11841] = 255;
assign img[11842] = 255;
assign img[11843] = 255;
assign img[11844] = 255;
assign img[11845] = 255;
assign img[11846] = 238;
assign img[11847] = 238;
assign img[11848] = 238;
assign img[11849] = 255;
assign img[11850] = 238;
assign img[11851] = 255;
assign img[11852] = 238;
assign img[11853] = 255;
assign img[11854] = 238;
assign img[11855] = 255;
assign img[11856] = 238;
assign img[11857] = 238;
assign img[11858] = 238;
assign img[11859] = 255;
assign img[11860] = 255;
assign img[11861] = 239;
assign img[11862] = 238;
assign img[11863] = 238;
assign img[11864] = 254;
assign img[11865] = 255;
assign img[11866] = 255;
assign img[11867] = 255;
assign img[11868] = 255;
assign img[11869] = 255;
assign img[11870] = 255;
assign img[11871] = 239;
assign img[11872] = 254;
assign img[11873] = 255;
assign img[11874] = 238;
assign img[11875] = 238;
assign img[11876] = 238;
assign img[11877] = 255;
assign img[11878] = 238;
assign img[11879] = 238;
assign img[11880] = 254;
assign img[11881] = 255;
assign img[11882] = 255;
assign img[11883] = 239;
assign img[11884] = 254;
assign img[11885] = 255;
assign img[11886] = 255;
assign img[11887] = 255;
assign img[11888] = 255;
assign img[11889] = 255;
assign img[11890] = 255;
assign img[11891] = 255;
assign img[11892] = 187;
assign img[11893] = 223;
assign img[11894] = 236;
assign img[11895] = 238;
assign img[11896] = 238;
assign img[11897] = 238;
assign img[11898] = 255;
assign img[11899] = 238;
assign img[11900] = 204;
assign img[11901] = 253;
assign img[11902] = 255;
assign img[11903] = 255;
assign img[11904] = 96;
assign img[11905] = 238;
assign img[11906] = 238;
assign img[11907] = 238;
assign img[11908] = 170;
assign img[11909] = 234;
assign img[11910] = 220;
assign img[11911] = 253;
assign img[11912] = 255;
assign img[11913] = 239;
assign img[11914] = 204;
assign img[11915] = 140;
assign img[11916] = 136;
assign img[11917] = 204;
assign img[11918] = 204;
assign img[11919] = 238;
assign img[11920] = 170;
assign img[11921] = 170;
assign img[11922] = 238;
assign img[11923] = 238;
assign img[11924] = 238;
assign img[11925] = 255;
assign img[11926] = 255;
assign img[11927] = 255;
assign img[11928] = 255;
assign img[11929] = 191;
assign img[11930] = 187;
assign img[11931] = 255;
assign img[11932] = 255;
assign img[11933] = 255;
assign img[11934] = 255;
assign img[11935] = 191;
assign img[11936] = 171;
assign img[11937] = 255;
assign img[11938] = 255;
assign img[11939] = 255;
assign img[11940] = 255;
assign img[11941] = 239;
assign img[11942] = 254;
assign img[11943] = 255;
assign img[11944] = 255;
assign img[11945] = 255;
assign img[11946] = 223;
assign img[11947] = 223;
assign img[11948] = 221;
assign img[11949] = 221;
assign img[11950] = 236;
assign img[11951] = 206;
assign img[11952] = 253;
assign img[11953] = 255;
assign img[11954] = 255;
assign img[11955] = 223;
assign img[11956] = 255;
assign img[11957] = 254;
assign img[11958] = 238;
assign img[11959] = 255;
assign img[11960] = 255;
assign img[11961] = 255;
assign img[11962] = 239;
assign img[11963] = 238;
assign img[11964] = 206;
assign img[11965] = 206;
assign img[11966] = 238;
assign img[11967] = 255;
assign img[11968] = 255;
assign img[11969] = 255;
assign img[11970] = 255;
assign img[11971] = 239;
assign img[11972] = 238;
assign img[11973] = 239;
assign img[11974] = 238;
assign img[11975] = 238;
assign img[11976] = 254;
assign img[11977] = 255;
assign img[11978] = 255;
assign img[11979] = 239;
assign img[11980] = 254;
assign img[11981] = 255;
assign img[11982] = 255;
assign img[11983] = 255;
assign img[11984] = 223;
assign img[11985] = 255;
assign img[11986] = 239;
assign img[11987] = 206;
assign img[11988] = 220;
assign img[11989] = 205;
assign img[11990] = 236;
assign img[11991] = 238;
assign img[11992] = 238;
assign img[11993] = 238;
assign img[11994] = 238;
assign img[11995] = 238;
assign img[11996] = 238;
assign img[11997] = 238;
assign img[11998] = 254;
assign img[11999] = 255;
assign img[12000] = 255;
assign img[12001] = 238;
assign img[12002] = 254;
assign img[12003] = 255;
assign img[12004] = 255;
assign img[12005] = 239;
assign img[12006] = 238;
assign img[12007] = 238;
assign img[12008] = 238;
assign img[12009] = 255;
assign img[12010] = 221;
assign img[12011] = 253;
assign img[12012] = 255;
assign img[12013] = 255;
assign img[12014] = 255;
assign img[12015] = 255;
assign img[12016] = 255;
assign img[12017] = 223;
assign img[12018] = 221;
assign img[12019] = 221;
assign img[12020] = 141;
assign img[12021] = 136;
assign img[12022] = 200;
assign img[12023] = 236;
assign img[12024] = 238;
assign img[12025] = 238;
assign img[12026] = 220;
assign img[12027] = 220;
assign img[12028] = 221;
assign img[12029] = 254;
assign img[12030] = 255;
assign img[12031] = 255;
assign img[12032] = 96;
assign img[12033] = 239;
assign img[12034] = 238;
assign img[12035] = 191;
assign img[12036] = 139;
assign img[12037] = 238;
assign img[12038] = 174;
assign img[12039] = 238;
assign img[12040] = 238;
assign img[12041] = 238;
assign img[12042] = 238;
assign img[12043] = 255;
assign img[12044] = 239;
assign img[12045] = 206;
assign img[12046] = 252;
assign img[12047] = 255;
assign img[12048] = 239;
assign img[12049] = 254;
assign img[12050] = 255;
assign img[12051] = 255;
assign img[12052] = 221;
assign img[12053] = 255;
assign img[12054] = 238;
assign img[12055] = 238;
assign img[12056] = 238;
assign img[12057] = 255;
assign img[12058] = 187;
assign img[12059] = 255;
assign img[12060] = 255;
assign img[12061] = 255;
assign img[12062] = 255;
assign img[12063] = 239;
assign img[12064] = 174;
assign img[12065] = 238;
assign img[12066] = 238;
assign img[12067] = 255;
assign img[12068] = 255;
assign img[12069] = 255;
assign img[12070] = 255;
assign img[12071] = 255;
assign img[12072] = 255;
assign img[12073] = 255;
assign img[12074] = 255;
assign img[12075] = 255;
assign img[12076] = 255;
assign img[12077] = 255;
assign img[12078] = 255;
assign img[12079] = 239;
assign img[12080] = 238;
assign img[12081] = 238;
assign img[12082] = 238;
assign img[12083] = 238;
assign img[12084] = 238;
assign img[12085] = 238;
assign img[12086] = 238;
assign img[12087] = 238;
assign img[12088] = 238;
assign img[12089] = 238;
assign img[12090] = 206;
assign img[12091] = 238;
assign img[12092] = 238;
assign img[12093] = 174;
assign img[12094] = 170;
assign img[12095] = 254;
assign img[12096] = 255;
assign img[12097] = 255;
assign img[12098] = 255;
assign img[12099] = 255;
assign img[12100] = 255;
assign img[12101] = 255;
assign img[12102] = 255;
assign img[12103] = 239;
assign img[12104] = 238;
assign img[12105] = 238;
assign img[12106] = 238;
assign img[12107] = 255;
assign img[12108] = 238;
assign img[12109] = 255;
assign img[12110] = 255;
assign img[12111] = 255;
assign img[12112] = 255;
assign img[12113] = 255;
assign img[12114] = 255;
assign img[12115] = 239;
assign img[12116] = 238;
assign img[12117] = 238;
assign img[12118] = 206;
assign img[12119] = 238;
assign img[12120] = 238;
assign img[12121] = 254;
assign img[12122] = 238;
assign img[12123] = 255;
assign img[12124] = 255;
assign img[12125] = 255;
assign img[12126] = 255;
assign img[12127] = 239;
assign img[12128] = 138;
assign img[12129] = 152;
assign img[12130] = 253;
assign img[12131] = 255;
assign img[12132] = 255;
assign img[12133] = 239;
assign img[12134] = 238;
assign img[12135] = 238;
assign img[12136] = 238;
assign img[12137] = 255;
assign img[12138] = 238;
assign img[12139] = 238;
assign img[12140] = 206;
assign img[12141] = 238;
assign img[12142] = 238;
assign img[12143] = 207;
assign img[12144] = 220;
assign img[12145] = 253;
assign img[12146] = 255;
assign img[12147] = 255;
assign img[12148] = 204;
assign img[12149] = 255;
assign img[12150] = 255;
assign img[12151] = 255;
assign img[12152] = 255;
assign img[12153] = 255;
assign img[12154] = 255;
assign img[12155] = 255;
assign img[12156] = 255;
assign img[12157] = 255;
assign img[12158] = 239;
assign img[12159] = 238;
assign img[12160] = 16;
assign img[12161] = 137;
assign img[12162] = 232;
assign img[12163] = 206;
assign img[12164] = 204;
assign img[12165] = 205;
assign img[12166] = 204;
assign img[12167] = 236;
assign img[12168] = 238;
assign img[12169] = 238;
assign img[12170] = 254;
assign img[12171] = 239;
assign img[12172] = 254;
assign img[12173] = 239;
assign img[12174] = 174;
assign img[12175] = 170;
assign img[12176] = 238;
assign img[12177] = 238;
assign img[12178] = 238;
assign img[12179] = 223;
assign img[12180] = 204;
assign img[12181] = 238;
assign img[12182] = 206;
assign img[12183] = 204;
assign img[12184] = 236;
assign img[12185] = 223;
assign img[12186] = 204;
assign img[12187] = 204;
assign img[12188] = 236;
assign img[12189] = 255;
assign img[12190] = 255;
assign img[12191] = 143;
assign img[12192] = 168;
assign img[12193] = 255;
assign img[12194] = 255;
assign img[12195] = 255;
assign img[12196] = 255;
assign img[12197] = 255;
assign img[12198] = 255;
assign img[12199] = 207;
assign img[12200] = 236;
assign img[12201] = 238;
assign img[12202] = 254;
assign img[12203] = 255;
assign img[12204] = 255;
assign img[12205] = 239;
assign img[12206] = 238;
assign img[12207] = 255;
assign img[12208] = 255;
assign img[12209] = 255;
assign img[12210] = 255;
assign img[12211] = 239;
assign img[12212] = 238;
assign img[12213] = 254;
assign img[12214] = 255;
assign img[12215] = 254;
assign img[12216] = 238;
assign img[12217] = 255;
assign img[12218] = 206;
assign img[12219] = 238;
assign img[12220] = 238;
assign img[12221] = 238;
assign img[12222] = 238;
assign img[12223] = 255;
assign img[12224] = 255;
assign img[12225] = 255;
assign img[12226] = 255;
assign img[12227] = 255;
assign img[12228] = 255;
assign img[12229] = 223;
assign img[12230] = 238;
assign img[12231] = 238;
assign img[12232] = 238;
assign img[12233] = 254;
assign img[12234] = 255;
assign img[12235] = 255;
assign img[12236] = 255;
assign img[12237] = 255;
assign img[12238] = 255;
assign img[12239] = 255;
assign img[12240] = 255;
assign img[12241] = 255;
assign img[12242] = 223;
assign img[12243] = 221;
assign img[12244] = 253;
assign img[12245] = 255;
assign img[12246] = 255;
assign img[12247] = 255;
assign img[12248] = 239;
assign img[12249] = 238;
assign img[12250] = 238;
assign img[12251] = 238;
assign img[12252] = 238;
assign img[12253] = 238;
assign img[12254] = 255;
assign img[12255] = 239;
assign img[12256] = 138;
assign img[12257] = 136;
assign img[12258] = 248;
assign img[12259] = 255;
assign img[12260] = 255;
assign img[12261] = 223;
assign img[12262] = 205;
assign img[12263] = 238;
assign img[12264] = 254;
assign img[12265] = 255;
assign img[12266] = 255;
assign img[12267] = 255;
assign img[12268] = 238;
assign img[12269] = 238;
assign img[12270] = 238;
assign img[12271] = 238;
assign img[12272] = 238;
assign img[12273] = 174;
assign img[12274] = 234;
assign img[12275] = 206;
assign img[12276] = 204;
assign img[12277] = 253;
assign img[12278] = 255;
assign img[12279] = 255;
assign img[12280] = 255;
assign img[12281] = 255;
assign img[12282] = 238;
assign img[12283] = 220;
assign img[12284] = 221;
assign img[12285] = 253;
assign img[12286] = 223;
assign img[12287] = 221;
assign img[12288] = 96;
assign img[12289] = 238;
assign img[12290] = 254;
assign img[12291] = 223;
assign img[12292] = 239;
assign img[12293] = 238;
assign img[12294] = 190;
assign img[12295] = 187;
assign img[12296] = 234;
assign img[12297] = 238;
assign img[12298] = 255;
assign img[12299] = 255;
assign img[12300] = 221;
assign img[12301] = 221;
assign img[12302] = 221;
assign img[12303] = 255;
assign img[12304] = 255;
assign img[12305] = 255;
assign img[12306] = 238;
assign img[12307] = 238;
assign img[12308] = 238;
assign img[12309] = 238;
assign img[12310] = 222;
assign img[12311] = 255;
assign img[12312] = 255;
assign img[12313] = 239;
assign img[12314] = 204;
assign img[12315] = 236;
assign img[12316] = 238;
assign img[12317] = 255;
assign img[12318] = 255;
assign img[12319] = 223;
assign img[12320] = 255;
assign img[12321] = 255;
assign img[12322] = 255;
assign img[12323] = 255;
assign img[12324] = 255;
assign img[12325] = 239;
assign img[12326] = 238;
assign img[12327] = 238;
assign img[12328] = 238;
assign img[12329] = 238;
assign img[12330] = 238;
assign img[12331] = 238;
assign img[12332] = 238;
assign img[12333] = 238;
assign img[12334] = 238;
assign img[12335] = 255;
assign img[12336] = 255;
assign img[12337] = 255;
assign img[12338] = 255;
assign img[12339] = 255;
assign img[12340] = 255;
assign img[12341] = 255;
assign img[12342] = 255;
assign img[12343] = 223;
assign img[12344] = 255;
assign img[12345] = 255;
assign img[12346] = 223;
assign img[12347] = 255;
assign img[12348] = 255;
assign img[12349] = 255;
assign img[12350] = 255;
assign img[12351] = 255;
assign img[12352] = 255;
assign img[12353] = 255;
assign img[12354] = 223;
assign img[12355] = 255;
assign img[12356] = 255;
assign img[12357] = 239;
assign img[12358] = 254;
assign img[12359] = 255;
assign img[12360] = 223;
assign img[12361] = 255;
assign img[12362] = 255;
assign img[12363] = 255;
assign img[12364] = 255;
assign img[12365] = 239;
assign img[12366] = 238;
assign img[12367] = 255;
assign img[12368] = 255;
assign img[12369] = 255;
assign img[12370] = 223;
assign img[12371] = 255;
assign img[12372] = 238;
assign img[12373] = 255;
assign img[12374] = 255;
assign img[12375] = 255;
assign img[12376] = 255;
assign img[12377] = 255;
assign img[12378] = 255;
assign img[12379] = 255;
assign img[12380] = 255;
assign img[12381] = 255;
assign img[12382] = 255;
assign img[12383] = 191;
assign img[12384] = 139;
assign img[12385] = 170;
assign img[12386] = 250;
assign img[12387] = 255;
assign img[12388] = 255;
assign img[12389] = 255;
assign img[12390] = 255;
assign img[12391] = 255;
assign img[12392] = 255;
assign img[12393] = 255;
assign img[12394] = 255;
assign img[12395] = 207;
assign img[12396] = 220;
assign img[12397] = 253;
assign img[12398] = 255;
assign img[12399] = 255;
assign img[12400] = 239;
assign img[12401] = 238;
assign img[12402] = 186;
assign img[12403] = 239;
assign img[12404] = 238;
assign img[12405] = 238;
assign img[12406] = 238;
assign img[12407] = 238;
assign img[12408] = 238;
assign img[12409] = 238;
assign img[12410] = 238;
assign img[12411] = 238;
assign img[12412] = 254;
assign img[12413] = 255;
assign img[12414] = 255;
assign img[12415] = 255;
assign img[12416] = 80;
assign img[12417] = 85;
assign img[12418] = 117;
assign img[12419] = 223;
assign img[12420] = 221;
assign img[12421] = 253;
assign img[12422] = 255;
assign img[12423] = 255;
assign img[12424] = 255;
assign img[12425] = 255;
assign img[12426] = 255;
assign img[12427] = 255;
assign img[12428] = 255;
assign img[12429] = 255;
assign img[12430] = 187;
assign img[12431] = 219;
assign img[12432] = 221;
assign img[12433] = 254;
assign img[12434] = 238;
assign img[12435] = 255;
assign img[12436] = 223;
assign img[12437] = 255;
assign img[12438] = 255;
assign img[12439] = 255;
assign img[12440] = 255;
assign img[12441] = 191;
assign img[12442] = 187;
assign img[12443] = 255;
assign img[12444] = 255;
assign img[12445] = 255;
assign img[12446] = 255;
assign img[12447] = 191;
assign img[12448] = 205;
assign img[12449] = 253;
assign img[12450] = 255;
assign img[12451] = 255;
assign img[12452] = 255;
assign img[12453] = 207;
assign img[12454] = 252;
assign img[12455] = 255;
assign img[12456] = 255;
assign img[12457] = 255;
assign img[12458] = 239;
assign img[12459] = 254;
assign img[12460] = 255;
assign img[12461] = 255;
assign img[12462] = 255;
assign img[12463] = 255;
assign img[12464] = 255;
assign img[12465] = 255;
assign img[12466] = 255;
assign img[12467] = 255;
assign img[12468] = 238;
assign img[12469] = 238;
assign img[12470] = 238;
assign img[12471] = 254;
assign img[12472] = 238;
assign img[12473] = 255;
assign img[12474] = 206;
assign img[12475] = 255;
assign img[12476] = 254;
assign img[12477] = 255;
assign img[12478] = 238;
assign img[12479] = 255;
assign img[12480] = 255;
assign img[12481] = 255;
assign img[12482] = 239;
assign img[12483] = 238;
assign img[12484] = 238;
assign img[12485] = 255;
assign img[12486] = 255;
assign img[12487] = 255;
assign img[12488] = 255;
assign img[12489] = 255;
assign img[12490] = 255;
assign img[12491] = 255;
assign img[12492] = 239;
assign img[12493] = 238;
assign img[12494] = 238;
assign img[12495] = 238;
assign img[12496] = 238;
assign img[12497] = 238;
assign img[12498] = 238;
assign img[12499] = 255;
assign img[12500] = 238;
assign img[12501] = 255;
assign img[12502] = 238;
assign img[12503] = 238;
assign img[12504] = 222;
assign img[12505] = 255;
assign img[12506] = 207;
assign img[12507] = 253;
assign img[12508] = 255;
assign img[12509] = 255;
assign img[12510] = 255;
assign img[12511] = 223;
assign img[12512] = 204;
assign img[12513] = 254;
assign img[12514] = 238;
assign img[12515] = 255;
assign img[12516] = 238;
assign img[12517] = 223;
assign img[12518] = 255;
assign img[12519] = 223;
assign img[12520] = 255;
assign img[12521] = 255;
assign img[12522] = 255;
assign img[12523] = 255;
assign img[12524] = 255;
assign img[12525] = 255;
assign img[12526] = 255;
assign img[12527] = 239;
assign img[12528] = 238;
assign img[12529] = 255;
assign img[12530] = 238;
assign img[12531] = 255;
assign img[12532] = 221;
assign img[12533] = 255;
assign img[12534] = 255;
assign img[12535] = 255;
assign img[12536] = 255;
assign img[12537] = 239;
assign img[12538] = 254;
assign img[12539] = 207;
assign img[12540] = 204;
assign img[12541] = 236;
assign img[12542] = 223;
assign img[12543] = 221;
assign img[12544] = 96;
assign img[12545] = 207;
assign img[12546] = 253;
assign img[12547] = 191;
assign img[12548] = 155;
assign img[12549] = 153;
assign img[12550] = 249;
assign img[12551] = 255;
assign img[12552] = 255;
assign img[12553] = 255;
assign img[12554] = 255;
assign img[12555] = 255;
assign img[12556] = 255;
assign img[12557] = 255;
assign img[12558] = 205;
assign img[12559] = 204;
assign img[12560] = 204;
assign img[12561] = 238;
assign img[12562] = 254;
assign img[12563] = 255;
assign img[12564] = 255;
assign img[12565] = 255;
assign img[12566] = 255;
assign img[12567] = 255;
assign img[12568] = 255;
assign img[12569] = 255;
assign img[12570] = 255;
assign img[12571] = 255;
assign img[12572] = 239;
assign img[12573] = 254;
assign img[12574] = 255;
assign img[12575] = 255;
assign img[12576] = 187;
assign img[12577] = 255;
assign img[12578] = 255;
assign img[12579] = 255;
assign img[12580] = 223;
assign img[12581] = 221;
assign img[12582] = 253;
assign img[12583] = 255;
assign img[12584] = 255;
assign img[12585] = 255;
assign img[12586] = 255;
assign img[12587] = 255;
assign img[12588] = 255;
assign img[12589] = 255;
assign img[12590] = 255;
assign img[12591] = 255;
assign img[12592] = 255;
assign img[12593] = 255;
assign img[12594] = 255;
assign img[12595] = 255;
assign img[12596] = 255;
assign img[12597] = 255;
assign img[12598] = 255;
assign img[12599] = 255;
assign img[12600] = 255;
assign img[12601] = 255;
assign img[12602] = 255;
assign img[12603] = 255;
assign img[12604] = 255;
assign img[12605] = 255;
assign img[12606] = 255;
assign img[12607] = 255;
assign img[12608] = 255;
assign img[12609] = 255;
assign img[12610] = 239;
assign img[12611] = 238;
assign img[12612] = 238;
assign img[12613] = 255;
assign img[12614] = 206;
assign img[12615] = 238;
assign img[12616] = 238;
assign img[12617] = 255;
assign img[12618] = 255;
assign img[12619] = 255;
assign img[12620] = 255;
assign img[12621] = 255;
assign img[12622] = 255;
assign img[12623] = 255;
assign img[12624] = 239;
assign img[12625] = 238;
assign img[12626] = 238;
assign img[12627] = 238;
assign img[12628] = 238;
assign img[12629] = 255;
assign img[12630] = 255;
assign img[12631] = 255;
assign img[12632] = 255;
assign img[12633] = 255;
assign img[12634] = 255;
assign img[12635] = 239;
assign img[12636] = 254;
assign img[12637] = 255;
assign img[12638] = 255;
assign img[12639] = 255;
assign img[12640] = 255;
assign img[12641] = 255;
assign img[12642] = 255;
assign img[12643] = 255;
assign img[12644] = 255;
assign img[12645] = 239;
assign img[12646] = 238;
assign img[12647] = 238;
assign img[12648] = 238;
assign img[12649] = 255;
assign img[12650] = 255;
assign img[12651] = 239;
assign img[12652] = 238;
assign img[12653] = 238;
assign img[12654] = 238;
assign img[12655] = 255;
assign img[12656] = 255;
assign img[12657] = 255;
assign img[12658] = 238;
assign img[12659] = 255;
assign img[12660] = 255;
assign img[12661] = 255;
assign img[12662] = 255;
assign img[12663] = 255;
assign img[12664] = 255;
assign img[12665] = 255;
assign img[12666] = 255;
assign img[12667] = 223;
assign img[12668] = 221;
assign img[12669] = 255;
assign img[12670] = 239;
assign img[12671] = 238;
assign img[12672] = 96;
assign img[12673] = 206;
assign img[12674] = 236;
assign img[12675] = 238;
assign img[12676] = 255;
assign img[12677] = 255;
assign img[12678] = 175;
assign img[12679] = 186;
assign img[12680] = 251;
assign img[12681] = 255;
assign img[12682] = 255;
assign img[12683] = 239;
assign img[12684] = 238;
assign img[12685] = 238;
assign img[12686] = 238;
assign img[12687] = 238;
assign img[12688] = 254;
assign img[12689] = 255;
assign img[12690] = 255;
assign img[12691] = 239;
assign img[12692] = 170;
assign img[12693] = 238;
assign img[12694] = 238;
assign img[12695] = 238;
assign img[12696] = 238;
assign img[12697] = 223;
assign img[12698] = 221;
assign img[12699] = 221;
assign img[12700] = 221;
assign img[12701] = 255;
assign img[12702] = 207;
assign img[12703] = 205;
assign img[12704] = 204;
assign img[12705] = 252;
assign img[12706] = 255;
assign img[12707] = 255;
assign img[12708] = 238;
assign img[12709] = 254;
assign img[12710] = 238;
assign img[12711] = 255;
assign img[12712] = 220;
assign img[12713] = 252;
assign img[12714] = 206;
assign img[12715] = 238;
assign img[12716] = 238;
assign img[12717] = 238;
assign img[12718] = 206;
assign img[12719] = 204;
assign img[12720] = 236;
assign img[12721] = 238;
assign img[12722] = 238;
assign img[12723] = 238;
assign img[12724] = 255;
assign img[12725] = 255;
assign img[12726] = 238;
assign img[12727] = 238;
assign img[12728] = 204;
assign img[12729] = 238;
assign img[12730] = 238;
assign img[12731] = 238;
assign img[12732] = 238;
assign img[12733] = 206;
assign img[12734] = 238;
assign img[12735] = 238;
assign img[12736] = 238;
assign img[12737] = 238;
assign img[12738] = 206;
assign img[12739] = 254;
assign img[12740] = 238;
assign img[12741] = 255;
assign img[12742] = 254;
assign img[12743] = 255;
assign img[12744] = 255;
assign img[12745] = 238;
assign img[12746] = 238;
assign img[12747] = 238;
assign img[12748] = 238;
assign img[12749] = 206;
assign img[12750] = 238;
assign img[12751] = 238;
assign img[12752] = 238;
assign img[12753] = 255;
assign img[12754] = 255;
assign img[12755] = 255;
assign img[12756] = 238;
assign img[12757] = 255;
assign img[12758] = 238;
assign img[12759] = 206;
assign img[12760] = 220;
assign img[12761] = 253;
assign img[12762] = 255;
assign img[12763] = 239;
assign img[12764] = 170;
assign img[12765] = 238;
assign img[12766] = 254;
assign img[12767] = 255;
assign img[12768] = 204;
assign img[12769] = 204;
assign img[12770] = 252;
assign img[12771] = 239;
assign img[12772] = 254;
assign img[12773] = 223;
assign img[12774] = 205;
assign img[12775] = 236;
assign img[12776] = 238;
assign img[12777] = 239;
assign img[12778] = 238;
assign img[12779] = 239;
assign img[12780] = 254;
assign img[12781] = 254;
assign img[12782] = 254;
assign img[12783] = 191;
assign img[12784] = 154;
assign img[12785] = 153;
assign img[12786] = 137;
assign img[12787] = 204;
assign img[12788] = 204;
assign img[12789] = 238;
assign img[12790] = 238;
assign img[12791] = 238;
assign img[12792] = 238;
assign img[12793] = 191;
assign img[12794] = 238;
assign img[12795] = 238;
assign img[12796] = 254;
assign img[12797] = 255;
assign img[12798] = 223;
assign img[12799] = 255;
assign img[12800] = 96;
assign img[12801] = 255;
assign img[12802] = 255;
assign img[12803] = 255;
assign img[12804] = 155;
assign img[12805] = 223;
assign img[12806] = 221;
assign img[12807] = 255;
assign img[12808] = 255;
assign img[12809] = 255;
assign img[12810] = 255;
assign img[12811] = 239;
assign img[12812] = 238;
assign img[12813] = 238;
assign img[12814] = 238;
assign img[12815] = 174;
assign img[12816] = 170;
assign img[12817] = 238;
assign img[12818] = 254;
assign img[12819] = 191;
assign img[12820] = 187;
assign img[12821] = 255;
assign img[12822] = 255;
assign img[12823] = 255;
assign img[12824] = 223;
assign img[12825] = 221;
assign img[12826] = 204;
assign img[12827] = 236;
assign img[12828] = 238;
assign img[12829] = 255;
assign img[12830] = 255;
assign img[12831] = 223;
assign img[12832] = 253;
assign img[12833] = 255;
assign img[12834] = 255;
assign img[12835] = 255;
assign img[12836] = 255;
assign img[12837] = 239;
assign img[12838] = 238;
assign img[12839] = 238;
assign img[12840] = 254;
assign img[12841] = 255;
assign img[12842] = 255;
assign img[12843] = 255;
assign img[12844] = 255;
assign img[12845] = 255;
assign img[12846] = 255;
assign img[12847] = 223;
assign img[12848] = 255;
assign img[12849] = 255;
assign img[12850] = 255;
assign img[12851] = 255;
assign img[12852] = 255;
assign img[12853] = 255;
assign img[12854] = 255;
assign img[12855] = 255;
assign img[12856] = 255;
assign img[12857] = 255;
assign img[12858] = 255;
assign img[12859] = 255;
assign img[12860] = 255;
assign img[12861] = 255;
assign img[12862] = 239;
assign img[12863] = 255;
assign img[12864] = 255;
assign img[12865] = 223;
assign img[12866] = 221;
assign img[12867] = 255;
assign img[12868] = 255;
assign img[12869] = 255;
assign img[12870] = 255;
assign img[12871] = 255;
assign img[12872] = 255;
assign img[12873] = 255;
assign img[12874] = 255;
assign img[12875] = 255;
assign img[12876] = 255;
assign img[12877] = 255;
assign img[12878] = 255;
assign img[12879] = 255;
assign img[12880] = 223;
assign img[12881] = 255;
assign img[12882] = 223;
assign img[12883] = 255;
assign img[12884] = 255;
assign img[12885] = 255;
assign img[12886] = 255;
assign img[12887] = 255;
assign img[12888] = 221;
assign img[12889] = 255;
assign img[12890] = 255;
assign img[12891] = 255;
assign img[12892] = 255;
assign img[12893] = 255;
assign img[12894] = 255;
assign img[12895] = 223;
assign img[12896] = 253;
assign img[12897] = 255;
assign img[12898] = 255;
assign img[12899] = 255;
assign img[12900] = 255;
assign img[12901] = 255;
assign img[12902] = 239;
assign img[12903] = 206;
assign img[12904] = 236;
assign img[12905] = 238;
assign img[12906] = 238;
assign img[12907] = 238;
assign img[12908] = 254;
assign img[12909] = 255;
assign img[12910] = 255;
assign img[12911] = 255;
assign img[12912] = 175;
assign img[12913] = 138;
assign img[12914] = 216;
assign img[12915] = 221;
assign img[12916] = 221;
assign img[12917] = 253;
assign img[12918] = 255;
assign img[12919] = 255;
assign img[12920] = 255;
assign img[12921] = 255;
assign img[12922] = 187;
assign img[12923] = 155;
assign img[12924] = 221;
assign img[12925] = 255;
assign img[12926] = 223;
assign img[12927] = 253;
assign img[12928] = 64;
assign img[12929] = 228;
assign img[12930] = 206;
assign img[12931] = 204;
assign img[12932] = 220;
assign img[12933] = 221;
assign img[12934] = 221;
assign img[12935] = 255;
assign img[12936] = 255;
assign img[12937] = 255;
assign img[12938] = 255;
assign img[12939] = 255;
assign img[12940] = 187;
assign img[12941] = 255;
assign img[12942] = 205;
assign img[12943] = 254;
assign img[12944] = 205;
assign img[12945] = 204;
assign img[12946] = 238;
assign img[12947] = 238;
assign img[12948] = 206;
assign img[12949] = 221;
assign img[12950] = 189;
assign img[12951] = 255;
assign img[12952] = 255;
assign img[12953] = 239;
assign img[12954] = 238;
assign img[12955] = 238;
assign img[12956] = 238;
assign img[12957] = 255;
assign img[12958] = 255;
assign img[12959] = 223;
assign img[12960] = 236;
assign img[12961] = 238;
assign img[12962] = 238;
assign img[12963] = 255;
assign img[12964] = 255;
assign img[12965] = 255;
assign img[12966] = 255;
assign img[12967] = 255;
assign img[12968] = 255;
assign img[12969] = 255;
assign img[12970] = 255;
assign img[12971] = 255;
assign img[12972] = 238;
assign img[12973] = 238;
assign img[12974] = 238;
assign img[12975] = 255;
assign img[12976] = 254;
assign img[12977] = 254;
assign img[12978] = 254;
assign img[12979] = 255;
assign img[12980] = 255;
assign img[12981] = 255;
assign img[12982] = 255;
assign img[12983] = 255;
assign img[12984] = 255;
assign img[12985] = 255;
assign img[12986] = 223;
assign img[12987] = 255;
assign img[12988] = 255;
assign img[12989] = 223;
assign img[12990] = 204;
assign img[12991] = 255;
assign img[12992] = 255;
assign img[12993] = 255;
assign img[12994] = 239;
assign img[12995] = 238;
assign img[12996] = 238;
assign img[12997] = 255;
assign img[12998] = 255;
assign img[12999] = 255;
assign img[13000] = 255;
assign img[13001] = 255;
assign img[13002] = 255;
assign img[13003] = 255;
assign img[13004] = 255;
assign img[13005] = 255;
assign img[13006] = 255;
assign img[13007] = 255;
assign img[13008] = 255;
assign img[13009] = 255;
assign img[13010] = 255;
assign img[13011] = 255;
assign img[13012] = 239;
assign img[13013] = 238;
assign img[13014] = 238;
assign img[13015] = 238;
assign img[13016] = 238;
assign img[13017] = 255;
assign img[13018] = 255;
assign img[13019] = 255;
assign img[13020] = 255;
assign img[13021] = 255;
assign img[13022] = 254;
assign img[13023] = 191;
assign img[13024] = 139;
assign img[13025] = 238;
assign img[13026] = 254;
assign img[13027] = 255;
assign img[13028] = 255;
assign img[13029] = 191;
assign img[13030] = 187;
assign img[13031] = 171;
assign img[13032] = 234;
assign img[13033] = 238;
assign img[13034] = 170;
assign img[13035] = 238;
assign img[13036] = 220;
assign img[13037] = 255;
assign img[13038] = 255;
assign img[13039] = 239;
assign img[13040] = 238;
assign img[13041] = 238;
assign img[13042] = 238;
assign img[13043] = 255;
assign img[13044] = 255;
assign img[13045] = 255;
assign img[13046] = 255;
assign img[13047] = 255;
assign img[13048] = 255;
assign img[13049] = 255;
assign img[13050] = 187;
assign img[13051] = 255;
assign img[13052] = 221;
assign img[13053] = 205;
assign img[13054] = 236;
assign img[13055] = 255;
assign img[13056] = 96;
assign img[13057] = 239;
assign img[13058] = 254;
assign img[13059] = 254;
assign img[13060] = 238;
assign img[13061] = 254;
assign img[13062] = 255;
assign img[13063] = 255;
assign img[13064] = 255;
assign img[13065] = 255;
assign img[13066] = 239;
assign img[13067] = 206;
assign img[13068] = 236;
assign img[13069] = 238;
assign img[13070] = 238;
assign img[13071] = 255;
assign img[13072] = 239;
assign img[13073] = 255;
assign img[13074] = 255;
assign img[13075] = 239;
assign img[13076] = 254;
assign img[13077] = 255;
assign img[13078] = 239;
assign img[13079] = 238;
assign img[13080] = 238;
assign img[13081] = 206;
assign img[13082] = 204;
assign img[13083] = 238;
assign img[13084] = 238;
assign img[13085] = 255;
assign img[13086] = 255;
assign img[13087] = 255;
assign img[13088] = 255;
assign img[13089] = 255;
assign img[13090] = 239;
assign img[13091] = 238;
assign img[13092] = 206;
assign img[13093] = 238;
assign img[13094] = 254;
assign img[13095] = 255;
assign img[13096] = 255;
assign img[13097] = 255;
assign img[13098] = 255;
assign img[13099] = 239;
assign img[13100] = 238;
assign img[13101] = 238;
assign img[13102] = 238;
assign img[13103] = 238;
assign img[13104] = 255;
assign img[13105] = 255;
assign img[13106] = 255;
assign img[13107] = 239;
assign img[13108] = 206;
assign img[13109] = 255;
assign img[13110] = 255;
assign img[13111] = 255;
assign img[13112] = 255;
assign img[13113] = 255;
assign img[13114] = 207;
assign img[13115] = 255;
assign img[13116] = 255;
assign img[13117] = 255;
assign img[13118] = 238;
assign img[13119] = 255;
assign img[13120] = 255;
assign img[13121] = 255;
assign img[13122] = 239;
assign img[13123] = 238;
assign img[13124] = 254;
assign img[13125] = 223;
assign img[13126] = 238;
assign img[13127] = 238;
assign img[13128] = 238;
assign img[13129] = 238;
assign img[13130] = 255;
assign img[13131] = 239;
assign img[13132] = 204;
assign img[13133] = 221;
assign img[13134] = 191;
assign img[13135] = 255;
assign img[13136] = 255;
assign img[13137] = 255;
assign img[13138] = 255;
assign img[13139] = 255;
assign img[13140] = 239;
assign img[13141] = 238;
assign img[13142] = 238;
assign img[13143] = 238;
assign img[13144] = 254;
assign img[13145] = 255;
assign img[13146] = 239;
assign img[13147] = 255;
assign img[13148] = 255;
assign img[13149] = 255;
assign img[13150] = 255;
assign img[13151] = 255;
assign img[13152] = 255;
assign img[13153] = 255;
assign img[13154] = 255;
assign img[13155] = 255;
assign img[13156] = 255;
assign img[13157] = 255;
assign img[13158] = 223;
assign img[13159] = 255;
assign img[13160] = 255;
assign img[13161] = 255;
assign img[13162] = 238;
assign img[13163] = 238;
assign img[13164] = 255;
assign img[13165] = 255;
assign img[13166] = 206;
assign img[13167] = 255;
assign img[13168] = 255;
assign img[13169] = 255;
assign img[13170] = 255;
assign img[13171] = 255;
assign img[13172] = 206;
assign img[13173] = 223;
assign img[13174] = 255;
assign img[13175] = 255;
assign img[13176] = 255;
assign img[13177] = 255;
assign img[13178] = 155;
assign img[13179] = 187;
assign img[13180] = 238;
assign img[13181] = 238;
assign img[13182] = 238;
assign img[13183] = 238;
assign img[13184] = 0;
assign img[13185] = 136;
assign img[13186] = 232;
assign img[13187] = 206;
assign img[13188] = 236;
assign img[13189] = 206;
assign img[13190] = 252;
assign img[13191] = 255;
assign img[13192] = 255;
assign img[13193] = 255;
assign img[13194] = 255;
assign img[13195] = 239;
assign img[13196] = 238;
assign img[13197] = 238;
assign img[13198] = 238;
assign img[13199] = 223;
assign img[13200] = 236;
assign img[13201] = 238;
assign img[13202] = 238;
assign img[13203] = 238;
assign img[13204] = 238;
assign img[13205] = 238;
assign img[13206] = 254;
assign img[13207] = 255;
assign img[13208] = 239;
assign img[13209] = 190;
assign img[13210] = 187;
assign img[13211] = 255;
assign img[13212] = 255;
assign img[13213] = 255;
assign img[13214] = 223;
assign img[13215] = 205;
assign img[13216] = 236;
assign img[13217] = 238;
assign img[13218] = 238;
assign img[13219] = 255;
assign img[13220] = 238;
assign img[13221] = 255;
assign img[13222] = 255;
assign img[13223] = 255;
assign img[13224] = 238;
assign img[13225] = 255;
assign img[13226] = 223;
assign img[13227] = 205;
assign img[13228] = 204;
assign img[13229] = 206;
assign img[13230] = 238;
assign img[13231] = 238;
assign img[13232] = 238;
assign img[13233] = 238;
assign img[13234] = 254;
assign img[13235] = 255;
assign img[13236] = 255;
assign img[13237] = 255;
assign img[13238] = 255;
assign img[13239] = 255;
assign img[13240] = 255;
assign img[13241] = 255;
assign img[13242] = 238;
assign img[13243] = 255;
assign img[13244] = 254;
assign img[13245] = 255;
assign img[13246] = 255;
assign img[13247] = 255;
assign img[13248] = 255;
assign img[13249] = 255;
assign img[13250] = 255;
assign img[13251] = 255;
assign img[13252] = 254;
assign img[13253] = 255;
assign img[13254] = 255;
assign img[13255] = 255;
assign img[13256] = 255;
assign img[13257] = 255;
assign img[13258] = 255;
assign img[13259] = 255;
assign img[13260] = 255;
assign img[13261] = 255;
assign img[13262] = 255;
assign img[13263] = 255;
assign img[13264] = 255;
assign img[13265] = 255;
assign img[13266] = 255;
assign img[13267] = 255;
assign img[13268] = 255;
assign img[13269] = 223;
assign img[13270] = 255;
assign img[13271] = 255;
assign img[13272] = 255;
assign img[13273] = 255;
assign img[13274] = 255;
assign img[13275] = 255;
assign img[13276] = 239;
assign img[13277] = 238;
assign img[13278] = 238;
assign img[13279] = 255;
assign img[13280] = 255;
assign img[13281] = 239;
assign img[13282] = 254;
assign img[13283] = 255;
assign img[13284] = 255;
assign img[13285] = 239;
assign img[13286] = 174;
assign img[13287] = 171;
assign img[13288] = 234;
assign img[13289] = 238;
assign img[13290] = 238;
assign img[13291] = 255;
assign img[13292] = 255;
assign img[13293] = 255;
assign img[13294] = 255;
assign img[13295] = 255;
assign img[13296] = 223;
assign img[13297] = 221;
assign img[13298] = 253;
assign img[13299] = 255;
assign img[13300] = 221;
assign img[13301] = 253;
assign img[13302] = 255;
assign img[13303] = 255;
assign img[13304] = 221;
assign img[13305] = 255;
assign img[13306] = 223;
assign img[13307] = 239;
assign img[13308] = 206;
assign img[13309] = 238;
assign img[13310] = 174;
assign img[13311] = 155;
assign img[13312] = 96;
assign img[13313] = 238;
assign img[13314] = 204;
assign img[13315] = 220;
assign img[13316] = 221;
assign img[13317] = 221;
assign img[13318] = 221;
assign img[13319] = 221;
assign img[13320] = 221;
assign img[13321] = 253;
assign img[13322] = 255;
assign img[13323] = 221;
assign img[13324] = 253;
assign img[13325] = 255;
assign img[13326] = 255;
assign img[13327] = 255;
assign img[13328] = 223;
assign img[13329] = 221;
assign img[13330] = 221;
assign img[13331] = 191;
assign img[13332] = 187;
assign img[13333] = 255;
assign img[13334] = 254;
assign img[13335] = 255;
assign img[13336] = 238;
assign img[13337] = 174;
assign img[13338] = 170;
assign img[13339] = 234;
assign img[13340] = 238;
assign img[13341] = 255;
assign img[13342] = 255;
assign img[13343] = 255;
assign img[13344] = 255;
assign img[13345] = 255;
assign img[13346] = 255;
assign img[13347] = 255;
assign img[13348] = 255;
assign img[13349] = 255;
assign img[13350] = 255;
assign img[13351] = 239;
assign img[13352] = 238;
assign img[13353] = 238;
assign img[13354] = 206;
assign img[13355] = 204;
assign img[13356] = 236;
assign img[13357] = 255;
assign img[13358] = 255;
assign img[13359] = 239;
assign img[13360] = 238;
assign img[13361] = 238;
assign img[13362] = 238;
assign img[13363] = 238;
assign img[13364] = 238;
assign img[13365] = 238;
assign img[13366] = 238;
assign img[13367] = 254;
assign img[13368] = 238;
assign img[13369] = 255;
assign img[13370] = 255;
assign img[13371] = 255;
assign img[13372] = 255;
assign img[13373] = 255;
assign img[13374] = 255;
assign img[13375] = 255;
assign img[13376] = 255;
assign img[13377] = 255;
assign img[13378] = 206;
assign img[13379] = 238;
assign img[13380] = 238;
assign img[13381] = 255;
assign img[13382] = 254;
assign img[13383] = 255;
assign img[13384] = 255;
assign img[13385] = 255;
assign img[13386] = 255;
assign img[13387] = 255;
assign img[13388] = 255;
assign img[13389] = 255;
assign img[13390] = 255;
assign img[13391] = 255;
assign img[13392] = 239;
assign img[13393] = 238;
assign img[13394] = 206;
assign img[13395] = 238;
assign img[13396] = 238;
assign img[13397] = 255;
assign img[13398] = 255;
assign img[13399] = 255;
assign img[13400] = 255;
assign img[13401] = 255;
assign img[13402] = 223;
assign img[13403] = 221;
assign img[13404] = 253;
assign img[13405] = 223;
assign img[13406] = 253;
assign img[13407] = 239;
assign img[13408] = 238;
assign img[13409] = 238;
assign img[13410] = 254;
assign img[13411] = 255;
assign img[13412] = 255;
assign img[13413] = 174;
assign img[13414] = 170;
assign img[13415] = 234;
assign img[13416] = 238;
assign img[13417] = 255;
assign img[13418] = 255;
assign img[13419] = 239;
assign img[13420] = 204;
assign img[13421] = 238;
assign img[13422] = 238;
assign img[13423] = 238;
assign img[13424] = 238;
assign img[13425] = 238;
assign img[13426] = 238;
assign img[13427] = 238;
assign img[13428] = 206;
assign img[13429] = 204;
assign img[13430] = 236;
assign img[13431] = 255;
assign img[13432] = 204;
assign img[13433] = 238;
assign img[13434] = 238;
assign img[13435] = 238;
assign img[13436] = 204;
assign img[13437] = 205;
assign img[13438] = 221;
assign img[13439] = 255;
assign img[13440] = 0;
assign img[13441] = 0;
assign img[13442] = 96;
assign img[13443] = 238;
assign img[13444] = 238;
assign img[13445] = 254;
assign img[13446] = 223;
assign img[13447] = 255;
assign img[13448] = 255;
assign img[13449] = 255;
assign img[13450] = 170;
assign img[13451] = 238;
assign img[13452] = 254;
assign img[13453] = 255;
assign img[13454] = 238;
assign img[13455] = 254;
assign img[13456] = 221;
assign img[13457] = 221;
assign img[13458] = 253;
assign img[13459] = 255;
assign img[13460] = 239;
assign img[13461] = 238;
assign img[13462] = 238;
assign img[13463] = 254;
assign img[13464] = 255;
assign img[13465] = 174;
assign img[13466] = 170;
assign img[13467] = 234;
assign img[13468] = 254;
assign img[13469] = 255;
assign img[13470] = 255;
assign img[13471] = 239;
assign img[13472] = 238;
assign img[13473] = 238;
assign img[13474] = 238;
assign img[13475] = 238;
assign img[13476] = 254;
assign img[13477] = 239;
assign img[13478] = 238;
assign img[13479] = 238;
assign img[13480] = 238;
assign img[13481] = 238;
assign img[13482] = 238;
assign img[13483] = 190;
assign img[13484] = 187;
assign img[13485] = 255;
assign img[13486] = 255;
assign img[13487] = 239;
assign img[13488] = 238;
assign img[13489] = 238;
assign img[13490] = 238;
assign img[13491] = 255;
assign img[13492] = 255;
assign img[13493] = 255;
assign img[13494] = 255;
assign img[13495] = 255;
assign img[13496] = 223;
assign img[13497] = 221;
assign img[13498] = 237;
assign img[13499] = 238;
assign img[13500] = 238;
assign img[13501] = 207;
assign img[13502] = 236;
assign img[13503] = 238;
assign img[13504] = 238;
assign img[13505] = 255;
assign img[13506] = 238;
assign img[13507] = 238;
assign img[13508] = 238;
assign img[13509] = 255;
assign img[13510] = 238;
assign img[13511] = 223;
assign img[13512] = 205;
assign img[13513] = 255;
assign img[13514] = 255;
assign img[13515] = 255;
assign img[13516] = 253;
assign img[13517] = 255;
assign img[13518] = 255;
assign img[13519] = 255;
assign img[13520] = 255;
assign img[13521] = 255;
assign img[13522] = 255;
assign img[13523] = 255;
assign img[13524] = 223;
assign img[13525] = 191;
assign img[13526] = 234;
assign img[13527] = 238;
assign img[13528] = 238;
assign img[13529] = 254;
assign img[13530] = 255;
assign img[13531] = 255;
assign img[13532] = 254;
assign img[13533] = 255;
assign img[13534] = 254;
assign img[13535] = 223;
assign img[13536] = 236;
assign img[13537] = 238;
assign img[13538] = 254;
assign img[13539] = 255;
assign img[13540] = 255;
assign img[13541] = 255;
assign img[13542] = 191;
assign img[13543] = 255;
assign img[13544] = 255;
assign img[13545] = 255;
assign img[13546] = 238;
assign img[13547] = 238;
assign img[13548] = 254;
assign img[13549] = 255;
assign img[13550] = 255;
assign img[13551] = 255;
assign img[13552] = 238;
assign img[13553] = 255;
assign img[13554] = 238;
assign img[13555] = 238;
assign img[13556] = 238;
assign img[13557] = 238;
assign img[13558] = 254;
assign img[13559] = 239;
assign img[13560] = 238;
assign img[13561] = 191;
assign img[13562] = 187;
assign img[13563] = 171;
assign img[13564] = 234;
assign img[13565] = 238;
assign img[13566] = 238;
assign img[13567] = 191;
assign img[13568] = 96;
assign img[13569] = 238;
assign img[13570] = 254;
assign img[13571] = 223;
assign img[13572] = 207;
assign img[13573] = 222;
assign img[13574] = 255;
assign img[13575] = 255;
assign img[13576] = 255;
assign img[13577] = 255;
assign img[13578] = 239;
assign img[13579] = 238;
assign img[13580] = 238;
assign img[13581] = 238;
assign img[13582] = 238;
assign img[13583] = 238;
assign img[13584] = 170;
assign img[13585] = 238;
assign img[13586] = 238;
assign img[13587] = 254;
assign img[13588] = 255;
assign img[13589] = 255;
assign img[13590] = 206;
assign img[13591] = 238;
assign img[13592] = 222;
assign img[13593] = 205;
assign img[13594] = 204;
assign img[13595] = 238;
assign img[13596] = 238;
assign img[13597] = 255;
assign img[13598] = 255;
assign img[13599] = 255;
assign img[13600] = 204;
assign img[13601] = 238;
assign img[13602] = 238;
assign img[13603] = 255;
assign img[13604] = 255;
assign img[13605] = 255;
assign img[13606] = 255;
assign img[13607] = 255;
assign img[13608] = 238;
assign img[13609] = 254;
assign img[13610] = 254;
assign img[13611] = 255;
assign img[13612] = 255;
assign img[13613] = 255;
assign img[13614] = 238;
assign img[13615] = 238;
assign img[13616] = 255;
assign img[13617] = 255;
assign img[13618] = 255;
assign img[13619] = 223;
assign img[13620] = 236;
assign img[13621] = 238;
assign img[13622] = 238;
assign img[13623] = 255;
assign img[13624] = 238;
assign img[13625] = 255;
assign img[13626] = 255;
assign img[13627] = 255;
assign img[13628] = 255;
assign img[13629] = 255;
assign img[13630] = 255;
assign img[13631] = 255;
assign img[13632] = 255;
assign img[13633] = 255;
assign img[13634] = 255;
assign img[13635] = 255;
assign img[13636] = 255;
assign img[13637] = 255;
assign img[13638] = 255;
assign img[13639] = 255;
assign img[13640] = 255;
assign img[13641] = 255;
assign img[13642] = 255;
assign img[13643] = 255;
assign img[13644] = 238;
assign img[13645] = 254;
assign img[13646] = 255;
assign img[13647] = 255;
assign img[13648] = 255;
assign img[13649] = 255;
assign img[13650] = 239;
assign img[13651] = 238;
assign img[13652] = 238;
assign img[13653] = 238;
assign img[13654] = 238;
assign img[13655] = 238;
assign img[13656] = 238;
assign img[13657] = 238;
assign img[13658] = 238;
assign img[13659] = 238;
assign img[13660] = 254;
assign img[13661] = 255;
assign img[13662] = 255;
assign img[13663] = 175;
assign img[13664] = 206;
assign img[13665] = 204;
assign img[13666] = 252;
assign img[13667] = 255;
assign img[13668] = 255;
assign img[13669] = 255;
assign img[13670] = 223;
assign img[13671] = 221;
assign img[13672] = 253;
assign img[13673] = 255;
assign img[13674] = 238;
assign img[13675] = 238;
assign img[13676] = 255;
assign img[13677] = 255;
assign img[13678] = 255;
assign img[13679] = 223;
assign img[13680] = 253;
assign img[13681] = 255;
assign img[13682] = 255;
assign img[13683] = 255;
assign img[13684] = 255;
assign img[13685] = 255;
assign img[13686] = 238;
assign img[13687] = 238;
assign img[13688] = 238;
assign img[13689] = 255;
assign img[13690] = 170;
assign img[13691] = 138;
assign img[13692] = 220;
assign img[13693] = 253;
assign img[13694] = 255;
assign img[13695] = 255;
assign img[13696] = 0;
assign img[13697] = 152;
assign img[13698] = 249;
assign img[13699] = 223;
assign img[13700] = 221;
assign img[13701] = 253;
assign img[13702] = 159;
assign img[13703] = 255;
assign img[13704] = 255;
assign img[13705] = 255;
assign img[13706] = 255;
assign img[13707] = 255;
assign img[13708] = 221;
assign img[13709] = 191;
assign img[13710] = 187;
assign img[13711] = 187;
assign img[13712] = 251;
assign img[13713] = 255;
assign img[13714] = 238;
assign img[13715] = 255;
assign img[13716] = 255;
assign img[13717] = 238;
assign img[13718] = 238;
assign img[13719] = 255;
assign img[13720] = 238;
assign img[13721] = 238;
assign img[13722] = 254;
assign img[13723] = 255;
assign img[13724] = 255;
assign img[13725] = 255;
assign img[13726] = 238;
assign img[13727] = 190;
assign img[13728] = 251;
assign img[13729] = 255;
assign img[13730] = 254;
assign img[13731] = 255;
assign img[13732] = 254;
assign img[13733] = 238;
assign img[13734] = 254;
assign img[13735] = 255;
assign img[13736] = 238;
assign img[13737] = 238;
assign img[13738] = 238;
assign img[13739] = 255;
assign img[13740] = 238;
assign img[13741] = 238;
assign img[13742] = 238;
assign img[13743] = 238;
assign img[13744] = 254;
assign img[13745] = 239;
assign img[13746] = 238;
assign img[13747] = 238;
assign img[13748] = 238;
assign img[13749] = 255;
assign img[13750] = 255;
assign img[13751] = 255;
assign img[13752] = 255;
assign img[13753] = 255;
assign img[13754] = 255;
assign img[13755] = 255;
assign img[13756] = 255;
assign img[13757] = 239;
assign img[13758] = 238;
assign img[13759] = 255;
assign img[13760] = 255;
assign img[13761] = 255;
assign img[13762] = 255;
assign img[13763] = 255;
assign img[13764] = 255;
assign img[13765] = 255;
assign img[13766] = 205;
assign img[13767] = 238;
assign img[13768] = 238;
assign img[13769] = 238;
assign img[13770] = 254;
assign img[13771] = 255;
assign img[13772] = 255;
assign img[13773] = 255;
assign img[13774] = 223;
assign img[13775] = 255;
assign img[13776] = 255;
assign img[13777] = 255;
assign img[13778] = 255;
assign img[13779] = 255;
assign img[13780] = 239;
assign img[13781] = 255;
assign img[13782] = 255;
assign img[13783] = 255;
assign img[13784] = 239;
assign img[13785] = 254;
assign img[13786] = 255;
assign img[13787] = 223;
assign img[13788] = 253;
assign img[13789] = 255;
assign img[13790] = 255;
assign img[13791] = 255;
assign img[13792] = 191;
assign img[13793] = 187;
assign img[13794] = 234;
assign img[13795] = 238;
assign img[13796] = 238;
assign img[13797] = 255;
assign img[13798] = 255;
assign img[13799] = 255;
assign img[13800] = 238;
assign img[13801] = 255;
assign img[13802] = 255;
assign img[13803] = 255;
assign img[13804] = 206;
assign img[13805] = 238;
assign img[13806] = 238;
assign img[13807] = 238;
assign img[13808] = 238;
assign img[13809] = 238;
assign img[13810] = 238;
assign img[13811] = 238;
assign img[13812] = 206;
assign img[13813] = 255;
assign img[13814] = 238;
assign img[13815] = 255;
assign img[13816] = 254;
assign img[13817] = 255;
assign img[13818] = 238;
assign img[13819] = 207;
assign img[13820] = 204;
assign img[13821] = 253;
assign img[13822] = 255;
assign img[13823] = 239;
assign img[13824] = 96;
assign img[13825] = 191;
assign img[13826] = 251;
assign img[13827] = 255;
assign img[13828] = 255;
assign img[13829] = 255;
assign img[13830] = 205;
assign img[13831] = 238;
assign img[13832] = 238;
assign img[13833] = 238;
assign img[13834] = 238;
assign img[13835] = 238;
assign img[13836] = 238;
assign img[13837] = 238;
assign img[13838] = 174;
assign img[13839] = 170;
assign img[13840] = 234;
assign img[13841] = 238;
assign img[13842] = 238;
assign img[13843] = 255;
assign img[13844] = 238;
assign img[13845] = 206;
assign img[13846] = 236;
assign img[13847] = 254;
assign img[13848] = 255;
assign img[13849] = 239;
assign img[13850] = 254;
assign img[13851] = 255;
assign img[13852] = 255;
assign img[13853] = 255;
assign img[13854] = 239;
assign img[13855] = 238;
assign img[13856] = 204;
assign img[13857] = 252;
assign img[13858] = 255;
assign img[13859] = 255;
assign img[13860] = 255;
assign img[13861] = 255;
assign img[13862] = 255;
assign img[13863] = 255;
assign img[13864] = 238;
assign img[13865] = 238;
assign img[13866] = 238;
assign img[13867] = 238;
assign img[13868] = 238;
assign img[13869] = 238;
assign img[13870] = 238;
assign img[13871] = 255;
assign img[13872] = 255;
assign img[13873] = 255;
assign img[13874] = 255;
assign img[13875] = 255;
assign img[13876] = 255;
assign img[13877] = 255;
assign img[13878] = 255;
assign img[13879] = 255;
assign img[13880] = 255;
assign img[13881] = 255;
assign img[13882] = 223;
assign img[13883] = 255;
assign img[13884] = 255;
assign img[13885] = 255;
assign img[13886] = 255;
assign img[13887] = 255;
assign img[13888] = 255;
assign img[13889] = 255;
assign img[13890] = 254;
assign img[13891] = 255;
assign img[13892] = 254;
assign img[13893] = 223;
assign img[13894] = 253;
assign img[13895] = 255;
assign img[13896] = 255;
assign img[13897] = 255;
assign img[13898] = 255;
assign img[13899] = 255;
assign img[13900] = 239;
assign img[13901] = 238;
assign img[13902] = 238;
assign img[13903] = 255;
assign img[13904] = 255;
assign img[13905] = 255;
assign img[13906] = 255;
assign img[13907] = 255;
assign img[13908] = 255;
assign img[13909] = 255;
assign img[13910] = 238;
assign img[13911] = 238;
assign img[13912] = 238;
assign img[13913] = 255;
assign img[13914] = 238;
assign img[13915] = 255;
assign img[13916] = 255;
assign img[13917] = 255;
assign img[13918] = 255;
assign img[13919] = 223;
assign img[13920] = 221;
assign img[13921] = 221;
assign img[13922] = 253;
assign img[13923] = 255;
assign img[13924] = 255;
assign img[13925] = 223;
assign img[13926] = 221;
assign img[13927] = 253;
assign img[13928] = 255;
assign img[13929] = 255;
assign img[13930] = 255;
assign img[13931] = 255;
assign img[13932] = 239;
assign img[13933] = 238;
assign img[13934] = 254;
assign img[13935] = 239;
assign img[13936] = 156;
assign img[13937] = 187;
assign img[13938] = 171;
assign img[13939] = 254;
assign img[13940] = 205;
assign img[13941] = 238;
assign img[13942] = 238;
assign img[13943] = 238;
assign img[13944] = 238;
assign img[13945] = 255;
assign img[13946] = 255;
assign img[13947] = 239;
assign img[13948] = 238;
assign img[13949] = 255;
assign img[13950] = 255;
assign img[13951] = 255;
assign img[13952] = 96;
assign img[13953] = 238;
assign img[13954] = 254;
assign img[13955] = 207;
assign img[13956] = 204;
assign img[13957] = 220;
assign img[13958] = 253;
assign img[13959] = 255;
assign img[13960] = 255;
assign img[13961] = 255;
assign img[13962] = 255;
assign img[13963] = 255;
assign img[13964] = 238;
assign img[13965] = 254;
assign img[13966] = 255;
assign img[13967] = 239;
assign img[13968] = 238;
assign img[13969] = 254;
assign img[13970] = 255;
assign img[13971] = 255;
assign img[13972] = 204;
assign img[13973] = 238;
assign img[13974] = 238;
assign img[13975] = 238;
assign img[13976] = 238;
assign img[13977] = 238;
assign img[13978] = 238;
assign img[13979] = 238;
assign img[13980] = 238;
assign img[13981] = 255;
assign img[13982] = 255;
assign img[13983] = 239;
assign img[13984] = 206;
assign img[13985] = 238;
assign img[13986] = 238;
assign img[13987] = 238;
assign img[13988] = 222;
assign img[13989] = 221;
assign img[13990] = 253;
assign img[13991] = 255;
assign img[13992] = 255;
assign img[13993] = 255;
assign img[13994] = 175;
assign img[13995] = 255;
assign img[13996] = 255;
assign img[13997] = 255;
assign img[13998] = 238;
assign img[13999] = 238;
assign img[14000] = 254;
assign img[14001] = 255;
assign img[14002] = 255;
assign img[14003] = 255;
assign img[14004] = 191;
assign img[14005] = 255;
assign img[14006] = 255;
assign img[14007] = 255;
assign img[14008] = 255;
assign img[14009] = 255;
assign img[14010] = 239;
assign img[14011] = 255;
assign img[14012] = 255;
assign img[14013] = 239;
assign img[14014] = 238;
assign img[14015] = 255;
assign img[14016] = 255;
assign img[14017] = 255;
assign img[14018] = 255;
assign img[14019] = 255;
assign img[14020] = 255;
assign img[14021] = 255;
assign img[14022] = 238;
assign img[14023] = 238;
assign img[14024] = 238;
assign img[14025] = 255;
assign img[14026] = 238;
assign img[14027] = 239;
assign img[14028] = 238;
assign img[14029] = 255;
assign img[14030] = 254;
assign img[14031] = 255;
assign img[14032] = 255;
assign img[14033] = 255;
assign img[14034] = 239;
assign img[14035] = 238;
assign img[14036] = 238;
assign img[14037] = 175;
assign img[14038] = 238;
assign img[14039] = 238;
assign img[14040] = 238;
assign img[14041] = 255;
assign img[14042] = 255;
assign img[14043] = 255;
assign img[14044] = 255;
assign img[14045] = 255;
assign img[14046] = 238;
assign img[14047] = 238;
assign img[14048] = 254;
assign img[14049] = 255;
assign img[14050] = 255;
assign img[14051] = 255;
assign img[14052] = 255;
assign img[14053] = 223;
assign img[14054] = 221;
assign img[14055] = 253;
assign img[14056] = 255;
assign img[14057] = 255;
assign img[14058] = 255;
assign img[14059] = 255;
assign img[14060] = 206;
assign img[14061] = 238;
assign img[14062] = 238;
assign img[14063] = 239;
assign img[14064] = 206;
assign img[14065] = 221;
assign img[14066] = 253;
assign img[14067] = 255;
assign img[14068] = 171;
assign img[14069] = 238;
assign img[14070] = 238;
assign img[14071] = 238;
assign img[14072] = 238;
assign img[14073] = 174;
assign img[14074] = 170;
assign img[14075] = 238;
assign img[14076] = 254;
assign img[14077] = 255;
assign img[14078] = 255;
assign img[14079] = 255;
assign img[14080] = 96;
assign img[14081] = 191;
assign img[14082] = 251;
assign img[14083] = 191;
assign img[14084] = 155;
assign img[14085] = 187;
assign img[14086] = 155;
assign img[14087] = 255;
assign img[14088] = 255;
assign img[14089] = 255;
assign img[14090] = 255;
assign img[14091] = 207;
assign img[14092] = 204;
assign img[14093] = 204;
assign img[14094] = 204;
assign img[14095] = 236;
assign img[14096] = 206;
assign img[14097] = 236;
assign img[14098] = 238;
assign img[14099] = 255;
assign img[14100] = 255;
assign img[14101] = 223;
assign img[14102] = 221;
assign img[14103] = 255;
assign img[14104] = 255;
assign img[14105] = 255;
assign img[14106] = 223;
assign img[14107] = 255;
assign img[14108] = 255;
assign img[14109] = 255;
assign img[14110] = 255;
assign img[14111] = 207;
assign img[14112] = 204;
assign img[14113] = 255;
assign img[14114] = 255;
assign img[14115] = 255;
assign img[14116] = 255;
assign img[14117] = 255;
assign img[14118] = 223;
assign img[14119] = 205;
assign img[14120] = 236;
assign img[14121] = 238;
assign img[14122] = 238;
assign img[14123] = 174;
assign img[14124] = 238;
assign img[14125] = 238;
assign img[14126] = 238;
assign img[14127] = 238;
assign img[14128] = 238;
assign img[14129] = 254;
assign img[14130] = 254;
assign img[14131] = 255;
assign img[14132] = 255;
assign img[14133] = 255;
assign img[14134] = 255;
assign img[14135] = 255;
assign img[14136] = 255;
assign img[14137] = 255;
assign img[14138] = 255;
assign img[14139] = 255;
assign img[14140] = 255;
assign img[14141] = 255;
assign img[14142] = 239;
assign img[14143] = 238;
assign img[14144] = 238;
assign img[14145] = 207;
assign img[14146] = 204;
assign img[14147] = 236;
assign img[14148] = 238;
assign img[14149] = 255;
assign img[14150] = 221;
assign img[14151] = 255;
assign img[14152] = 255;
assign img[14153] = 255;
assign img[14154] = 255;
assign img[14155] = 223;
assign img[14156] = 221;
assign img[14157] = 255;
assign img[14158] = 255;
assign img[14159] = 255;
assign img[14160] = 223;
assign img[14161] = 255;
assign img[14162] = 223;
assign img[14163] = 255;
assign img[14164] = 191;
assign img[14165] = 171;
assign img[14166] = 234;
assign img[14167] = 238;
assign img[14168] = 238;
assign img[14169] = 238;
assign img[14170] = 204;
assign img[14171] = 254;
assign img[14172] = 255;
assign img[14173] = 255;
assign img[14174] = 255;
assign img[14175] = 191;
assign img[14176] = 255;
assign img[14177] = 238;
assign img[14178] = 254;
assign img[14179] = 255;
assign img[14180] = 255;
assign img[14181] = 223;
assign img[14182] = 221;
assign img[14183] = 255;
assign img[14184] = 255;
assign img[14185] = 255;
assign img[14186] = 255;
assign img[14187] = 255;
assign img[14188] = 255;
assign img[14189] = 255;
assign img[14190] = 255;
assign img[14191] = 223;
assign img[14192] = 221;
assign img[14193] = 221;
assign img[14194] = 221;
assign img[14195] = 221;
assign img[14196] = 221;
assign img[14197] = 205;
assign img[14198] = 236;
assign img[14199] = 238;
assign img[14200] = 238;
assign img[14201] = 238;
assign img[14202] = 220;
assign img[14203] = 221;
assign img[14204] = 173;
assign img[14205] = 238;
assign img[14206] = 190;
assign img[14207] = 255;
assign img[14208] = 96;
assign img[14209] = 206;
assign img[14210] = 204;
assign img[14211] = 204;
assign img[14212] = 204;
assign img[14213] = 204;
assign img[14214] = 140;
assign img[14215] = 220;
assign img[14216] = 237;
assign img[14217] = 238;
assign img[14218] = 238;
assign img[14219] = 207;
assign img[14220] = 204;
assign img[14221] = 236;
assign img[14222] = 254;
assign img[14223] = 221;
assign img[14224] = 221;
assign img[14225] = 221;
assign img[14226] = 253;
assign img[14227] = 223;
assign img[14228] = 204;
assign img[14229] = 204;
assign img[14230] = 221;
assign img[14231] = 255;
assign img[14232] = 255;
assign img[14233] = 239;
assign img[14234] = 170;
assign img[14235] = 238;
assign img[14236] = 238;
assign img[14237] = 255;
assign img[14238] = 255;
assign img[14239] = 239;
assign img[14240] = 174;
assign img[14241] = 238;
assign img[14242] = 238;
assign img[14243] = 255;
assign img[14244] = 255;
assign img[14245] = 239;
assign img[14246] = 238;
assign img[14247] = 255;
assign img[14248] = 255;
assign img[14249] = 255;
assign img[14250] = 255;
assign img[14251] = 255;
assign img[14252] = 255;
assign img[14253] = 255;
assign img[14254] = 255;
assign img[14255] = 255;
assign img[14256] = 255;
assign img[14257] = 255;
assign img[14258] = 255;
assign img[14259] = 255;
assign img[14260] = 255;
assign img[14261] = 255;
assign img[14262] = 255;
assign img[14263] = 255;
assign img[14264] = 255;
assign img[14265] = 255;
assign img[14266] = 239;
assign img[14267] = 206;
assign img[14268] = 238;
assign img[14269] = 238;
assign img[14270] = 238;
assign img[14271] = 255;
assign img[14272] = 255;
assign img[14273] = 255;
assign img[14274] = 255;
assign img[14275] = 255;
assign img[14276] = 255;
assign img[14277] = 255;
assign img[14278] = 238;
assign img[14279] = 238;
assign img[14280] = 238;
assign img[14281] = 238;
assign img[14282] = 254;
assign img[14283] = 255;
assign img[14284] = 239;
assign img[14285] = 238;
assign img[14286] = 238;
assign img[14287] = 255;
assign img[14288] = 255;
assign img[14289] = 255;
assign img[14290] = 255;
assign img[14291] = 255;
assign img[14292] = 255;
assign img[14293] = 255;
assign img[14294] = 238;
assign img[14295] = 255;
assign img[14296] = 255;
assign img[14297] = 255;
assign img[14298] = 255;
assign img[14299] = 255;
assign img[14300] = 255;
assign img[14301] = 255;
assign img[14302] = 255;
assign img[14303] = 239;
assign img[14304] = 138;
assign img[14305] = 155;
assign img[14306] = 255;
assign img[14307] = 255;
assign img[14308] = 255;
assign img[14309] = 239;
assign img[14310] = 238;
assign img[14311] = 238;
assign img[14312] = 238;
assign img[14313] = 254;
assign img[14314] = 221;
assign img[14315] = 221;
assign img[14316] = 205;
assign img[14317] = 236;
assign img[14318] = 222;
assign img[14319] = 221;
assign img[14320] = 205;
assign img[14321] = 236;
assign img[14322] = 238;
assign img[14323] = 255;
assign img[14324] = 205;
assign img[14325] = 204;
assign img[14326] = 252;
assign img[14327] = 255;
assign img[14328] = 223;
assign img[14329] = 239;
assign img[14330] = 254;
assign img[14331] = 255;
assign img[14332] = 255;
assign img[14333] = 239;
assign img[14334] = 220;
assign img[14335] = 253;
assign img[14336] = 0;
assign img[14337] = 204;
assign img[14338] = 236;
assign img[14339] = 206;
assign img[14340] = 236;
assign img[14341] = 238;
assign img[14342] = 186;
assign img[14343] = 251;
assign img[14344] = 255;
assign img[14345] = 255;
assign img[14346] = 221;
assign img[14347] = 223;
assign img[14348] = 221;
assign img[14349] = 253;
assign img[14350] = 255;
assign img[14351] = 191;
assign img[14352] = 255;
assign img[14353] = 255;
assign img[14354] = 255;
assign img[14355] = 255;
assign img[14356] = 255;
assign img[14357] = 255;
assign img[14358] = 239;
assign img[14359] = 238;
assign img[14360] = 238;
assign img[14361] = 206;
assign img[14362] = 204;
assign img[14363] = 236;
assign img[14364] = 238;
assign img[14365] = 238;
assign img[14366] = 238;
assign img[14367] = 206;
assign img[14368] = 204;
assign img[14369] = 236;
assign img[14370] = 238;
assign img[14371] = 255;
assign img[14372] = 255;
assign img[14373] = 255;
assign img[14374] = 255;
assign img[14375] = 223;
assign img[14376] = 253;
assign img[14377] = 255;
assign img[14378] = 207;
assign img[14379] = 221;
assign img[14380] = 255;
assign img[14381] = 255;
assign img[14382] = 238;
assign img[14383] = 238;
assign img[14384] = 238;
assign img[14385] = 238;
assign img[14386] = 238;
assign img[14387] = 238;
assign img[14388] = 254;
assign img[14389] = 255;
assign img[14390] = 255;
assign img[14391] = 255;
assign img[14392] = 255;
assign img[14393] = 255;
assign img[14394] = 223;
assign img[14395] = 221;
assign img[14396] = 253;
assign img[14397] = 255;
assign img[14398] = 255;
assign img[14399] = 255;
assign img[14400] = 255;
assign img[14401] = 255;
assign img[14402] = 255;
assign img[14403] = 255;
assign img[14404] = 239;
assign img[14405] = 206;
assign img[14406] = 220;
assign img[14407] = 255;
assign img[14408] = 223;
assign img[14409] = 255;
assign img[14410] = 255;
assign img[14411] = 255;
assign img[14412] = 255;
assign img[14413] = 255;
assign img[14414] = 255;
assign img[14415] = 255;
assign img[14416] = 239;
assign img[14417] = 238;
assign img[14418] = 238;
assign img[14419] = 238;
assign img[14420] = 174;
assign img[14421] = 171;
assign img[14422] = 234;
assign img[14423] = 238;
assign img[14424] = 206;
assign img[14425] = 204;
assign img[14426] = 220;
assign img[14427] = 239;
assign img[14428] = 254;
assign img[14429] = 255;
assign img[14430] = 255;
assign img[14431] = 239;
assign img[14432] = 254;
assign img[14433] = 255;
assign img[14434] = 238;
assign img[14435] = 238;
assign img[14436] = 238;
assign img[14437] = 255;
assign img[14438] = 221;
assign img[14439] = 253;
assign img[14440] = 255;
assign img[14441] = 255;
assign img[14442] = 236;
assign img[14443] = 238;
assign img[14444] = 255;
assign img[14445] = 255;
assign img[14446] = 223;
assign img[14447] = 223;
assign img[14448] = 191;
assign img[14449] = 139;
assign img[14450] = 248;
assign img[14451] = 223;
assign img[14452] = 253;
assign img[14453] = 239;
assign img[14454] = 238;
assign img[14455] = 238;
assign img[14456] = 238;
assign img[14457] = 238;
assign img[14458] = 254;
assign img[14459] = 255;
assign img[14460] = 223;
assign img[14461] = 255;
assign img[14462] = 239;
assign img[14463] = 238;
assign img[14464] = 96;
assign img[14465] = 87;
assign img[14466] = 117;
assign img[14467] = 255;
assign img[14468] = 239;
assign img[14469] = 238;
assign img[14470] = 254;
assign img[14471] = 255;
assign img[14472] = 255;
assign img[14473] = 255;
assign img[14474] = 239;
assign img[14475] = 206;
assign img[14476] = 204;
assign img[14477] = 236;
assign img[14478] = 238;
assign img[14479] = 238;
assign img[14480] = 254;
assign img[14481] = 255;
assign img[14482] = 255;
assign img[14483] = 255;
assign img[14484] = 206;
assign img[14485] = 221;
assign img[14486] = 141;
assign img[14487] = 236;
assign img[14488] = 238;
assign img[14489] = 238;
assign img[14490] = 238;
assign img[14491] = 238;
assign img[14492] = 238;
assign img[14493] = 238;
assign img[14494] = 238;
assign img[14495] = 255;
assign img[14496] = 187;
assign img[14497] = 251;
assign img[14498] = 255;
assign img[14499] = 255;
assign img[14500] = 255;
assign img[14501] = 255;
assign img[14502] = 255;
assign img[14503] = 239;
assign img[14504] = 238;
assign img[14505] = 238;
assign img[14506] = 238;
assign img[14507] = 238;
assign img[14508] = 254;
assign img[14509] = 239;
assign img[14510] = 238;
assign img[14511] = 238;
assign img[14512] = 238;
assign img[14513] = 238;
assign img[14514] = 238;
assign img[14515] = 238;
assign img[14516] = 254;
assign img[14517] = 255;
assign img[14518] = 255;
assign img[14519] = 255;
assign img[14520] = 238;
assign img[14521] = 223;
assign img[14522] = 221;
assign img[14523] = 253;
assign img[14524] = 255;
assign img[14525] = 255;
assign img[14526] = 255;
assign img[14527] = 255;
assign img[14528] = 255;
assign img[14529] = 239;
assign img[14530] = 238;
assign img[14531] = 238;
assign img[14532] = 238;
assign img[14533] = 238;
assign img[14534] = 220;
assign img[14535] = 253;
assign img[14536] = 255;
assign img[14537] = 255;
assign img[14538] = 223;
assign img[14539] = 221;
assign img[14540] = 221;
assign img[14541] = 255;
assign img[14542] = 255;
assign img[14543] = 255;
assign img[14544] = 255;
assign img[14545] = 255;
assign img[14546] = 255;
assign img[14547] = 255;
assign img[14548] = 255;
assign img[14549] = 255;
assign img[14550] = 255;
assign img[14551] = 255;
assign img[14552] = 255;
assign img[14553] = 255;
assign img[14554] = 255;
assign img[14555] = 255;
assign img[14556] = 255;
assign img[14557] = 255;
assign img[14558] = 255;
assign img[14559] = 191;
assign img[14560] = 251;
assign img[14561] = 255;
assign img[14562] = 255;
assign img[14563] = 255;
assign img[14564] = 254;
assign img[14565] = 255;
assign img[14566] = 206;
assign img[14567] = 238;
assign img[14568] = 238;
assign img[14569] = 206;
assign img[14570] = 204;
assign img[14571] = 221;
assign img[14572] = 205;
assign img[14573] = 238;
assign img[14574] = 238;
assign img[14575] = 206;
assign img[14576] = 204;
assign img[14577] = 236;
assign img[14578] = 255;
assign img[14579] = 255;
assign img[14580] = 223;
assign img[14581] = 221;
assign img[14582] = 236;
assign img[14583] = 238;
assign img[14584] = 238;
assign img[14585] = 238;
assign img[14586] = 170;
assign img[14587] = 238;
assign img[14588] = 254;
assign img[14589] = 255;
assign img[14590] = 223;
assign img[14591] = 255;
assign img[14592] = 112;
assign img[14593] = 223;
assign img[14594] = 253;
assign img[14595] = 255;
assign img[14596] = 171;
assign img[14597] = 238;
assign img[14598] = 174;
assign img[14599] = 238;
assign img[14600] = 238;
assign img[14601] = 255;
assign img[14602] = 221;
assign img[14603] = 221;
assign img[14604] = 204;
assign img[14605] = 236;
assign img[14606] = 190;
assign img[14607] = 191;
assign img[14608] = 187;
assign img[14609] = 255;
assign img[14610] = 238;
assign img[14611] = 191;
assign img[14612] = 187;
assign img[14613] = 187;
assign img[14614] = 187;
assign img[14615] = 255;
assign img[14616] = 255;
assign img[14617] = 223;
assign img[14618] = 221;
assign img[14619] = 253;
assign img[14620] = 255;
assign img[14621] = 255;
assign img[14622] = 239;
assign img[14623] = 174;
assign img[14624] = 206;
assign img[14625] = 238;
assign img[14626] = 254;
assign img[14627] = 239;
assign img[14628] = 238;
assign img[14629] = 238;
assign img[14630] = 238;
assign img[14631] = 238;
assign img[14632] = 238;
assign img[14633] = 238;
assign img[14634] = 238;
assign img[14635] = 255;
assign img[14636] = 238;
assign img[14637] = 238;
assign img[14638] = 238;
assign img[14639] = 239;
assign img[14640] = 255;
assign img[14641] = 255;
assign img[14642] = 255;
assign img[14643] = 255;
assign img[14644] = 223;
assign img[14645] = 255;
assign img[14646] = 254;
assign img[14647] = 255;
assign img[14648] = 255;
assign img[14649] = 255;
assign img[14650] = 255;
assign img[14651] = 255;
assign img[14652] = 255;
assign img[14653] = 255;
assign img[14654] = 255;
assign img[14655] = 255;
assign img[14656] = 255;
assign img[14657] = 255;
assign img[14658] = 223;
assign img[14659] = 255;
assign img[14660] = 238;
assign img[14661] = 255;
assign img[14662] = 238;
assign img[14663] = 238;
assign img[14664] = 238;
assign img[14665] = 238;
assign img[14666] = 254;
assign img[14667] = 255;
assign img[14668] = 255;
assign img[14669] = 255;
assign img[14670] = 255;
assign img[14671] = 255;
assign img[14672] = 239;
assign img[14673] = 238;
assign img[14674] = 238;
assign img[14675] = 238;
assign img[14676] = 238;
assign img[14677] = 223;
assign img[14678] = 255;
assign img[14679] = 255;
assign img[14680] = 255;
assign img[14681] = 255;
assign img[14682] = 223;
assign img[14683] = 255;
assign img[14684] = 255;
assign img[14685] = 255;
assign img[14686] = 255;
assign img[14687] = 255;
assign img[14688] = 255;
assign img[14689] = 255;
assign img[14690] = 255;
assign img[14691] = 255;
assign img[14692] = 255;
assign img[14693] = 223;
assign img[14694] = 238;
assign img[14695] = 238;
assign img[14696] = 238;
assign img[14697] = 238;
assign img[14698] = 186;
assign img[14699] = 187;
assign img[14700] = 187;
assign img[14701] = 251;
assign img[14702] = 238;
assign img[14703] = 238;
assign img[14704] = 140;
assign img[14705] = 170;
assign img[14706] = 234;
assign img[14707] = 255;
assign img[14708] = 238;
assign img[14709] = 238;
assign img[14710] = 238;
assign img[14711] = 238;
assign img[14712] = 238;
assign img[14713] = 255;
assign img[14714] = 255;
assign img[14715] = 255;
assign img[14716] = 238;
assign img[14717] = 255;
assign img[14718] = 255;
assign img[14719] = 223;
assign img[14720] = 0;
assign img[14721] = 204;
assign img[14722] = 252;
assign img[14723] = 223;
assign img[14724] = 221;
assign img[14725] = 221;
assign img[14726] = 141;
assign img[14727] = 238;
assign img[14728] = 238;
assign img[14729] = 254;
assign img[14730] = 254;
assign img[14731] = 255;
assign img[14732] = 255;
assign img[14733] = 223;
assign img[14734] = 205;
assign img[14735] = 221;
assign img[14736] = 221;
assign img[14737] = 221;
assign img[14738] = 221;
assign img[14739] = 157;
assign img[14740] = 253;
assign img[14741] = 255;
assign img[14742] = 255;
assign img[14743] = 255;
assign img[14744] = 255;
assign img[14745] = 239;
assign img[14746] = 138;
assign img[14747] = 238;
assign img[14748] = 238;
assign img[14749] = 255;
assign img[14750] = 255;
assign img[14751] = 239;
assign img[14752] = 204;
assign img[14753] = 238;
assign img[14754] = 238;
assign img[14755] = 255;
assign img[14756] = 255;
assign img[14757] = 255;
assign img[14758] = 255;
assign img[14759] = 255;
assign img[14760] = 255;
assign img[14761] = 255;
assign img[14762] = 223;
assign img[14763] = 255;
assign img[14764] = 223;
assign img[14765] = 237;
assign img[14766] = 238;
assign img[14767] = 255;
assign img[14768] = 255;
assign img[14769] = 255;
assign img[14770] = 255;
assign img[14771] = 255;
assign img[14772] = 255;
assign img[14773] = 255;
assign img[14774] = 255;
assign img[14775] = 255;
assign img[14776] = 255;
assign img[14777] = 255;
assign img[14778] = 239;
assign img[14779] = 238;
assign img[14780] = 254;
assign img[14781] = 239;
assign img[14782] = 238;
assign img[14783] = 255;
assign img[14784] = 255;
assign img[14785] = 255;
assign img[14786] = 255;
assign img[14787] = 255;
assign img[14788] = 255;
assign img[14789] = 255;
assign img[14790] = 238;
assign img[14791] = 238;
assign img[14792] = 255;
assign img[14793] = 255;
assign img[14794] = 255;
assign img[14795] = 255;
assign img[14796] = 255;
assign img[14797] = 255;
assign img[14798] = 255;
assign img[14799] = 255;
assign img[14800] = 254;
assign img[14801] = 255;
assign img[14802] = 254;
assign img[14803] = 206;
assign img[14804] = 238;
assign img[14805] = 206;
assign img[14806] = 236;
assign img[14807] = 238;
assign img[14808] = 238;
assign img[14809] = 255;
assign img[14810] = 255;
assign img[14811] = 255;
assign img[14812] = 255;
assign img[14813] = 255;
assign img[14814] = 255;
assign img[14815] = 255;
assign img[14816] = 155;
assign img[14817] = 239;
assign img[14818] = 254;
assign img[14819] = 255;
assign img[14820] = 255;
assign img[14821] = 255;
assign img[14822] = 221;
assign img[14823] = 255;
assign img[14824] = 255;
assign img[14825] = 255;
assign img[14826] = 255;
assign img[14827] = 255;
assign img[14828] = 191;
assign img[14829] = 187;
assign img[14830] = 251;
assign img[14831] = 223;
assign img[14832] = 221;
assign img[14833] = 221;
assign img[14834] = 221;
assign img[14835] = 221;
assign img[14836] = 253;
assign img[14837] = 255;
assign img[14838] = 255;
assign img[14839] = 255;
assign img[14840] = 255;
assign img[14841] = 175;
assign img[14842] = 170;
assign img[14843] = 170;
assign img[14844] = 234;
assign img[14845] = 254;
assign img[14846] = 255;
assign img[14847] = 223;
assign img[14848] = 96;
assign img[14849] = 119;
assign img[14850] = 119;
assign img[14851] = 207;
assign img[14852] = 204;
assign img[14853] = 204;
assign img[14854] = 204;
assign img[14855] = 204;
assign img[14856] = 236;
assign img[14857] = 255;
assign img[14858] = 221;
assign img[14859] = 255;
assign img[14860] = 238;
assign img[14861] = 255;
assign img[14862] = 239;
assign img[14863] = 206;
assign img[14864] = 220;
assign img[14865] = 255;
assign img[14866] = 255;
assign img[14867] = 255;
assign img[14868] = 238;
assign img[14869] = 255;
assign img[14870] = 171;
assign img[14871] = 238;
assign img[14872] = 174;
assign img[14873] = 170;
assign img[14874] = 250;
assign img[14875] = 255;
assign img[14876] = 255;
assign img[14877] = 255;
assign img[14878] = 238;
assign img[14879] = 238;
assign img[14880] = 204;
assign img[14881] = 236;
assign img[14882] = 238;
assign img[14883] = 238;
assign img[14884] = 238;
assign img[14885] = 238;
assign img[14886] = 238;
assign img[14887] = 255;
assign img[14888] = 254;
assign img[14889] = 238;
assign img[14890] = 238;
assign img[14891] = 238;
assign img[14892] = 238;
assign img[14893] = 255;
assign img[14894] = 238;
assign img[14895] = 239;
assign img[14896] = 238;
assign img[14897] = 238;
assign img[14898] = 238;
assign img[14899] = 238;
assign img[14900] = 238;
assign img[14901] = 254;
assign img[14902] = 238;
assign img[14903] = 238;
assign img[14904] = 238;
assign img[14905] = 238;
assign img[14906] = 238;
assign img[14907] = 238;
assign img[14908] = 238;
assign img[14909] = 222;
assign img[14910] = 254;
assign img[14911] = 255;
assign img[14912] = 255;
assign img[14913] = 255;
assign img[14914] = 223;
assign img[14915] = 255;
assign img[14916] = 255;
assign img[14917] = 255;
assign img[14918] = 255;
assign img[14919] = 255;
assign img[14920] = 223;
assign img[14921] = 221;
assign img[14922] = 236;
assign img[14923] = 255;
assign img[14924] = 255;
assign img[14925] = 255;
assign img[14926] = 255;
assign img[14927] = 255;
assign img[14928] = 223;
assign img[14929] = 255;
assign img[14930] = 238;
assign img[14931] = 238;
assign img[14932] = 238;
assign img[14933] = 206;
assign img[14934] = 204;
assign img[14935] = 238;
assign img[14936] = 238;
assign img[14937] = 255;
assign img[14938] = 255;
assign img[14939] = 255;
assign img[14940] = 255;
assign img[14941] = 255;
assign img[14942] = 255;
assign img[14943] = 223;
assign img[14944] = 204;
assign img[14945] = 206;
assign img[14946] = 238;
assign img[14947] = 238;
assign img[14948] = 238;
assign img[14949] = 238;
assign img[14950] = 254;
assign img[14951] = 255;
assign img[14952] = 238;
assign img[14953] = 255;
assign img[14954] = 174;
assign img[14955] = 238;
assign img[14956] = 174;
assign img[14957] = 238;
assign img[14958] = 238;
assign img[14959] = 238;
assign img[14960] = 254;
assign img[14961] = 255;
assign img[14962] = 170;
assign img[14963] = 239;
assign img[14964] = 238;
assign img[14965] = 238;
assign img[14966] = 238;
assign img[14967] = 238;
assign img[14968] = 254;
assign img[14969] = 175;
assign img[14970] = 238;
assign img[14971] = 206;
assign img[14972] = 204;
assign img[14973] = 236;
assign img[14974] = 238;
assign img[14975] = 255;
assign img[14976] = 96;
assign img[14977] = 206;
assign img[14978] = 236;
assign img[14979] = 238;
assign img[14980] = 204;
assign img[14981] = 204;
assign img[14982] = 220;
assign img[14983] = 255;
assign img[14984] = 255;
assign img[14985] = 255;
assign img[14986] = 238;
assign img[14987] = 222;
assign img[14988] = 205;
assign img[14989] = 238;
assign img[14990] = 206;
assign img[14991] = 220;
assign img[14992] = 221;
assign img[14993] = 253;
assign img[14994] = 255;
assign img[14995] = 255;
assign img[14996] = 255;
assign img[14997] = 223;
assign img[14998] = 253;
assign img[14999] = 255;
assign img[15000] = 255;
assign img[15001] = 255;
assign img[15002] = 255;
assign img[15003] = 255;
assign img[15004] = 255;
assign img[15005] = 255;
assign img[15006] = 239;
assign img[15007] = 238;
assign img[15008] = 254;
assign img[15009] = 255;
assign img[15010] = 255;
assign img[15011] = 255;
assign img[15012] = 255;
assign img[15013] = 255;
assign img[15014] = 255;
assign img[15015] = 255;
assign img[15016] = 238;
assign img[15017] = 238;
assign img[15018] = 238;
assign img[15019] = 255;
assign img[15020] = 238;
assign img[15021] = 255;
assign img[15022] = 238;
assign img[15023] = 255;
assign img[15024] = 255;
assign img[15025] = 255;
assign img[15026] = 255;
assign img[15027] = 255;
assign img[15028] = 255;
assign img[15029] = 255;
assign img[15030] = 255;
assign img[15031] = 239;
assign img[15032] = 238;
assign img[15033] = 238;
assign img[15034] = 238;
assign img[15035] = 255;
assign img[15036] = 238;
assign img[15037] = 238;
assign img[15038] = 238;
assign img[15039] = 255;
assign img[15040] = 255;
assign img[15041] = 255;
assign img[15042] = 255;
assign img[15043] = 255;
assign img[15044] = 239;
assign img[15045] = 238;
assign img[15046] = 254;
assign img[15047] = 255;
assign img[15048] = 255;
assign img[15049] = 255;
assign img[15050] = 255;
assign img[15051] = 255;
assign img[15052] = 255;
assign img[15053] = 255;
assign img[15054] = 255;
assign img[15055] = 255;
assign img[15056] = 255;
assign img[15057] = 255;
assign img[15058] = 255;
assign img[15059] = 255;
assign img[15060] = 255;
assign img[15061] = 255;
assign img[15062] = 255;
assign img[15063] = 255;
assign img[15064] = 239;
assign img[15065] = 255;
assign img[15066] = 255;
assign img[15067] = 255;
assign img[15068] = 255;
assign img[15069] = 255;
assign img[15070] = 255;
assign img[15071] = 223;
assign img[15072] = 221;
assign img[15073] = 223;
assign img[15074] = 255;
assign img[15075] = 255;
assign img[15076] = 255;
assign img[15077] = 255;
assign img[15078] = 139;
assign img[15079] = 136;
assign img[15080] = 238;
assign img[15081] = 238;
assign img[15082] = 238;
assign img[15083] = 222;
assign img[15084] = 221;
assign img[15085] = 255;
assign img[15086] = 255;
assign img[15087] = 239;
assign img[15088] = 204;
assign img[15089] = 204;
assign img[15090] = 236;
assign img[15091] = 239;
assign img[15092] = 206;
assign img[15093] = 237;
assign img[15094] = 238;
assign img[15095] = 238;
assign img[15096] = 238;
assign img[15097] = 174;
assign img[15098] = 186;
assign img[15099] = 187;
assign img[15100] = 217;
assign img[15101] = 253;
assign img[15102] = 191;
assign img[15103] = 255;
assign img[15104] = 80;
assign img[15105] = 103;
assign img[15106] = 118;
assign img[15107] = 191;
assign img[15108] = 187;
assign img[15109] = 187;
assign img[15110] = 187;
assign img[15111] = 187;
assign img[15112] = 234;
assign img[15113] = 255;
assign img[15114] = 255;
assign img[15115] = 223;
assign img[15116] = 249;
assign img[15117] = 255;
assign img[15118] = 191;
assign img[15119] = 155;
assign img[15120] = 201;
assign img[15121] = 204;
assign img[15122] = 204;
assign img[15123] = 220;
assign img[15124] = 153;
assign img[15125] = 255;
assign img[15126] = 207;
assign img[15127] = 236;
assign img[15128] = 206;
assign img[15129] = 204;
assign img[15130] = 236;
assign img[15131] = 238;
assign img[15132] = 238;
assign img[15133] = 255;
assign img[15134] = 255;
assign img[15135] = 255;
assign img[15136] = 239;
assign img[15137] = 255;
assign img[15138] = 255;
assign img[15139] = 255;
assign img[15140] = 255;
assign img[15141] = 255;
assign img[15142] = 255;
assign img[15143] = 255;
assign img[15144] = 255;
assign img[15145] = 255;
assign img[15146] = 255;
assign img[15147] = 255;
assign img[15148] = 239;
assign img[15149] = 254;
assign img[15150] = 255;
assign img[15151] = 223;
assign img[15152] = 255;
assign img[15153] = 255;
assign img[15154] = 255;
assign img[15155] = 255;
assign img[15156] = 255;
assign img[15157] = 255;
assign img[15158] = 255;
assign img[15159] = 255;
assign img[15160] = 255;
assign img[15161] = 255;
assign img[15162] = 238;
assign img[15163] = 238;
assign img[15164] = 238;
assign img[15165] = 206;
assign img[15166] = 238;
assign img[15167] = 238;
assign img[15168] = 238;
assign img[15169] = 254;
assign img[15170] = 206;
assign img[15171] = 254;
assign img[15172] = 254;
assign img[15173] = 191;
assign img[15174] = 238;
assign img[15175] = 238;
assign img[15176] = 238;
assign img[15177] = 238;
assign img[15178] = 254;
assign img[15179] = 239;
assign img[15180] = 238;
assign img[15181] = 238;
assign img[15182] = 238;
assign img[15183] = 238;
assign img[15184] = 238;
assign img[15185] = 238;
assign img[15186] = 238;
assign img[15187] = 255;
assign img[15188] = 238;
assign img[15189] = 239;
assign img[15190] = 238;
assign img[15191] = 238;
assign img[15192] = 238;
assign img[15193] = 238;
assign img[15194] = 255;
assign img[15195] = 255;
assign img[15196] = 255;
assign img[15197] = 255;
assign img[15198] = 255;
assign img[15199] = 255;
assign img[15200] = 238;
assign img[15201] = 238;
assign img[15202] = 254;
assign img[15203] = 255;
assign img[15204] = 255;
assign img[15205] = 238;
assign img[15206] = 238;
assign img[15207] = 254;
assign img[15208] = 255;
assign img[15209] = 255;
assign img[15210] = 255;
assign img[15211] = 239;
assign img[15212] = 238;
assign img[15213] = 238;
assign img[15214] = 255;
assign img[15215] = 223;
assign img[15216] = 221;
assign img[15217] = 189;
assign img[15218] = 251;
assign img[15219] = 255;
assign img[15220] = 223;
assign img[15221] = 221;
assign img[15222] = 221;
assign img[15223] = 255;
assign img[15224] = 255;
assign img[15225] = 255;
assign img[15226] = 221;
assign img[15227] = 191;
assign img[15228] = 171;
assign img[15229] = 238;
assign img[15230] = 254;
assign img[15231] = 255;
assign img[15232] = 64;
assign img[15233] = 206;
assign img[15234] = 254;
assign img[15235] = 223;
assign img[15236] = 221;
assign img[15237] = 221;
assign img[15238] = 205;
assign img[15239] = 238;
assign img[15240] = 238;
assign img[15241] = 238;
assign img[15242] = 238;
assign img[15243] = 255;
assign img[15244] = 239;
assign img[15245] = 238;
assign img[15246] = 238;
assign img[15247] = 174;
assign img[15248] = 204;
assign img[15249] = 204;
assign img[15250] = 236;
assign img[15251] = 255;
assign img[15252] = 255;
assign img[15253] = 255;
assign img[15254] = 255;
assign img[15255] = 255;
assign img[15256] = 255;
assign img[15257] = 239;
assign img[15258] = 238;
assign img[15259] = 238;
assign img[15260] = 238;
assign img[15261] = 255;
assign img[15262] = 223;
assign img[15263] = 221;
assign img[15264] = 221;
assign img[15265] = 253;
assign img[15266] = 255;
assign img[15267] = 255;
assign img[15268] = 255;
assign img[15269] = 255;
assign img[15270] = 255;
assign img[15271] = 239;
assign img[15272] = 238;
assign img[15273] = 238;
assign img[15274] = 238;
assign img[15275] = 238;
assign img[15276] = 238;
assign img[15277] = 238;
assign img[15278] = 238;
assign img[15279] = 255;
assign img[15280] = 255;
assign img[15281] = 255;
assign img[15282] = 255;
assign img[15283] = 255;
assign img[15284] = 223;
assign img[15285] = 255;
assign img[15286] = 239;
assign img[15287] = 238;
assign img[15288] = 238;
assign img[15289] = 238;
assign img[15290] = 254;
assign img[15291] = 255;
assign img[15292] = 255;
assign img[15293] = 255;
assign img[15294] = 255;
assign img[15295] = 255;
assign img[15296] = 255;
assign img[15297] = 255;
assign img[15298] = 255;
assign img[15299] = 255;
assign img[15300] = 255;
assign img[15301] = 255;
assign img[15302] = 255;
assign img[15303] = 239;
assign img[15304] = 238;
assign img[15305] = 239;
assign img[15306] = 255;
assign img[15307] = 255;
assign img[15308] = 255;
assign img[15309] = 255;
assign img[15310] = 255;
assign img[15311] = 255;
assign img[15312] = 255;
assign img[15313] = 255;
assign img[15314] = 255;
assign img[15315] = 255;
assign img[15316] = 255;
assign img[15317] = 223;
assign img[15318] = 255;
assign img[15319] = 255;
assign img[15320] = 255;
assign img[15321] = 255;
assign img[15322] = 255;
assign img[15323] = 255;
assign img[15324] = 255;
assign img[15325] = 255;
assign img[15326] = 255;
assign img[15327] = 255;
assign img[15328] = 255;
assign img[15329] = 223;
assign img[15330] = 253;
assign img[15331] = 255;
assign img[15332] = 255;
assign img[15333] = 255;
assign img[15334] = 223;
assign img[15335] = 221;
assign img[15336] = 253;
assign img[15337] = 255;
assign img[15338] = 238;
assign img[15339] = 238;
assign img[15340] = 238;
assign img[15341] = 255;
assign img[15342] = 254;
assign img[15343] = 238;
assign img[15344] = 238;
assign img[15345] = 238;
assign img[15346] = 238;
assign img[15347] = 239;
assign img[15348] = 238;
assign img[15349] = 238;
assign img[15350] = 254;
assign img[15351] = 255;
assign img[15352] = 221;
assign img[15353] = 255;
assign img[15354] = 221;
assign img[15355] = 221;
assign img[15356] = 221;
assign img[15357] = 253;
assign img[15358] = 255;
assign img[15359] = 255;
assign img[15360] = 96;
assign img[15361] = 238;
assign img[15362] = 238;
assign img[15363] = 255;
assign img[15364] = 255;
assign img[15365] = 255;
assign img[15366] = 221;
assign img[15367] = 255;
assign img[15368] = 255;
assign img[15369] = 255;
assign img[15370] = 239;
assign img[15371] = 238;
assign img[15372] = 238;
assign img[15373] = 238;
assign img[15374] = 238;
assign img[15375] = 238;
assign img[15376] = 238;
assign img[15377] = 238;
assign img[15378] = 254;
assign img[15379] = 255;
assign img[15380] = 171;
assign img[15381] = 238;
assign img[15382] = 158;
assign img[15383] = 255;
assign img[15384] = 255;
assign img[15385] = 191;
assign img[15386] = 139;
assign img[15387] = 238;
assign img[15388] = 238;
assign img[15389] = 255;
assign img[15390] = 255;
assign img[15391] = 255;
assign img[15392] = 174;
assign img[15393] = 187;
assign img[15394] = 251;
assign img[15395] = 255;
assign img[15396] = 238;
assign img[15397] = 238;
assign img[15398] = 238;
assign img[15399] = 255;
assign img[15400] = 238;
assign img[15401] = 255;
assign img[15402] = 254;
assign img[15403] = 254;
assign img[15404] = 254;
assign img[15405] = 238;
assign img[15406] = 238;
assign img[15407] = 255;
assign img[15408] = 255;
assign img[15409] = 255;
assign img[15410] = 255;
assign img[15411] = 255;
assign img[15412] = 255;
assign img[15413] = 255;
assign img[15414] = 255;
assign img[15415] = 255;
assign img[15416] = 255;
assign img[15417] = 255;
assign img[15418] = 255;
assign img[15419] = 255;
assign img[15420] = 255;
assign img[15421] = 255;
assign img[15422] = 255;
assign img[15423] = 239;
assign img[15424] = 238;
assign img[15425] = 238;
assign img[15426] = 254;
assign img[15427] = 255;
assign img[15428] = 255;
assign img[15429] = 255;
assign img[15430] = 255;
assign img[15431] = 255;
assign img[15432] = 255;
assign img[15433] = 255;
assign img[15434] = 255;
assign img[15435] = 255;
assign img[15436] = 223;
assign img[15437] = 255;
assign img[15438] = 255;
assign img[15439] = 255;
assign img[15440] = 223;
assign img[15441] = 255;
assign img[15442] = 255;
assign img[15443] = 255;
assign img[15444] = 255;
assign img[15445] = 255;
assign img[15446] = 254;
assign img[15447] = 255;
assign img[15448] = 223;
assign img[15449] = 255;
assign img[15450] = 255;
assign img[15451] = 255;
assign img[15452] = 239;
assign img[15453] = 238;
assign img[15454] = 238;
assign img[15455] = 191;
assign img[15456] = 171;
assign img[15457] = 238;
assign img[15458] = 254;
assign img[15459] = 255;
assign img[15460] = 255;
assign img[15461] = 255;
assign img[15462] = 204;
assign img[15463] = 238;
assign img[15464] = 238;
assign img[15465] = 254;
assign img[15466] = 254;
assign img[15467] = 255;
assign img[15468] = 238;
assign img[15469] = 255;
assign img[15470] = 239;
assign img[15471] = 238;
assign img[15472] = 206;
assign img[15473] = 254;
assign img[15474] = 255;
assign img[15475] = 255;
assign img[15476] = 255;
assign img[15477] = 255;
assign img[15478] = 238;
assign img[15479] = 255;
assign img[15480] = 255;
assign img[15481] = 255;
assign img[15482] = 171;
assign img[15483] = 238;
assign img[15484] = 206;
assign img[15485] = 238;
assign img[15486] = 238;
assign img[15487] = 254;
assign img[15488] = 96;
assign img[15489] = 238;
assign img[15490] = 238;
assign img[15491] = 255;
assign img[15492] = 187;
assign img[15493] = 238;
assign img[15494] = 254;
assign img[15495] = 191;
assign img[15496] = 255;
assign img[15497] = 255;
assign img[15498] = 255;
assign img[15499] = 255;
assign img[15500] = 222;
assign img[15501] = 221;
assign img[15502] = 221;
assign img[15503] = 205;
assign img[15504] = 204;
assign img[15505] = 204;
assign img[15506] = 204;
assign img[15507] = 204;
assign img[15508] = 252;
assign img[15509] = 255;
assign img[15510] = 239;
assign img[15511] = 238;
assign img[15512] = 238;
assign img[15513] = 238;
assign img[15514] = 170;
assign img[15515] = 238;
assign img[15516] = 223;
assign img[15517] = 255;
assign img[15518] = 255;
assign img[15519] = 191;
assign img[15520] = 171;
assign img[15521] = 234;
assign img[15522] = 238;
assign img[15523] = 238;
assign img[15524] = 238;
assign img[15525] = 238;
assign img[15526] = 238;
assign img[15527] = 255;
assign img[15528] = 255;
assign img[15529] = 255;
assign img[15530] = 255;
assign img[15531] = 255;
assign img[15532] = 238;
assign img[15533] = 255;
assign img[15534] = 238;
assign img[15535] = 255;
assign img[15536] = 255;
assign img[15537] = 255;
assign img[15538] = 255;
assign img[15539] = 255;
assign img[15540] = 255;
assign img[15541] = 255;
assign img[15542] = 255;
assign img[15543] = 255;
assign img[15544] = 255;
assign img[15545] = 255;
assign img[15546] = 223;
assign img[15547] = 255;
assign img[15548] = 255;
assign img[15549] = 207;
assign img[15550] = 204;
assign img[15551] = 238;
assign img[15552] = 238;
assign img[15553] = 255;
assign img[15554] = 223;
assign img[15555] = 255;
assign img[15556] = 255;
assign img[15557] = 255;
assign img[15558] = 221;
assign img[15559] = 255;
assign img[15560] = 255;
assign img[15561] = 255;
assign img[15562] = 255;
assign img[15563] = 255;
assign img[15564] = 255;
assign img[15565] = 255;
assign img[15566] = 255;
assign img[15567] = 255;
assign img[15568] = 255;
assign img[15569] = 255;
assign img[15570] = 255;
assign img[15571] = 255;
assign img[15572] = 255;
assign img[15573] = 255;
assign img[15574] = 255;
assign img[15575] = 255;
assign img[15576] = 255;
assign img[15577] = 255;
assign img[15578] = 255;
assign img[15579] = 255;
assign img[15580] = 238;
assign img[15581] = 238;
assign img[15582] = 238;
assign img[15583] = 191;
assign img[15584] = 170;
assign img[15585] = 234;
assign img[15586] = 255;
assign img[15587] = 223;
assign img[15588] = 255;
assign img[15589] = 239;
assign img[15590] = 238;
assign img[15591] = 238;
assign img[15592] = 238;
assign img[15593] = 255;
assign img[15594] = 238;
assign img[15595] = 238;
assign img[15596] = 254;
assign img[15597] = 255;
assign img[15598] = 255;
assign img[15599] = 255;
assign img[15600] = 221;
assign img[15601] = 205;
assign img[15602] = 236;
assign img[15603] = 206;
assign img[15604] = 236;
assign img[15605] = 238;
assign img[15606] = 238;
assign img[15607] = 254;
assign img[15608] = 255;
assign img[15609] = 255;
assign img[15610] = 255;
assign img[15611] = 239;
assign img[15612] = 238;
assign img[15613] = 238;
assign img[15614] = 238;
assign img[15615] = 238;
assign img[15616] = 80;
assign img[15617] = 213;
assign img[15618] = 236;
assign img[15619] = 238;
assign img[15620] = 254;
assign img[15621] = 255;
assign img[15622] = 223;
assign img[15623] = 221;
assign img[15624] = 253;
assign img[15625] = 223;
assign img[15626] = 252;
assign img[15627] = 223;
assign img[15628] = 253;
assign img[15629] = 255;
assign img[15630] = 239;
assign img[15631] = 206;
assign img[15632] = 204;
assign img[15633] = 204;
assign img[15634] = 236;
assign img[15635] = 174;
assign img[15636] = 154;
assign img[15637] = 205;
assign img[15638] = 236;
assign img[15639] = 238;
assign img[15640] = 238;
assign img[15641] = 191;
assign img[15642] = 187;
assign img[15643] = 255;
assign img[15644] = 255;
assign img[15645] = 255;
assign img[15646] = 255;
assign img[15647] = 255;
assign img[15648] = 255;
assign img[15649] = 255;
assign img[15650] = 255;
assign img[15651] = 255;
assign img[15652] = 255;
assign img[15653] = 255;
assign img[15654] = 255;
assign img[15655] = 239;
assign img[15656] = 238;
assign img[15657] = 238;
assign img[15658] = 238;
assign img[15659] = 238;
assign img[15660] = 238;
assign img[15661] = 238;
assign img[15662] = 238;
assign img[15663] = 255;
assign img[15664] = 255;
assign img[15665] = 255;
assign img[15666] = 255;
assign img[15667] = 255;
assign img[15668] = 255;
assign img[15669] = 255;
assign img[15670] = 255;
assign img[15671] = 255;
assign img[15672] = 255;
assign img[15673] = 255;
assign img[15674] = 255;
assign img[15675] = 255;
assign img[15676] = 255;
assign img[15677] = 255;
assign img[15678] = 255;
assign img[15679] = 255;
assign img[15680] = 255;
assign img[15681] = 255;
assign img[15682] = 255;
assign img[15683] = 255;
assign img[15684] = 255;
assign img[15685] = 255;
assign img[15686] = 255;
assign img[15687] = 255;
assign img[15688] = 239;
assign img[15689] = 238;
assign img[15690] = 254;
assign img[15691] = 239;
assign img[15692] = 238;
assign img[15693] = 238;
assign img[15694] = 238;
assign img[15695] = 255;
assign img[15696] = 255;
assign img[15697] = 255;
assign img[15698] = 255;
assign img[15699] = 255;
assign img[15700] = 239;
assign img[15701] = 239;
assign img[15702] = 238;
assign img[15703] = 238;
assign img[15704] = 174;
assign img[15705] = 238;
assign img[15706] = 238;
assign img[15707] = 255;
assign img[15708] = 255;
assign img[15709] = 255;
assign img[15710] = 255;
assign img[15711] = 255;
assign img[15712] = 238;
assign img[15713] = 255;
assign img[15714] = 255;
assign img[15715] = 255;
assign img[15716] = 255;
assign img[15717] = 255;
assign img[15718] = 255;
assign img[15719] = 254;
assign img[15720] = 254;
assign img[15721] = 255;
assign img[15722] = 255;
assign img[15723] = 255;
assign img[15724] = 255;
assign img[15725] = 255;
assign img[15726] = 255;
assign img[15727] = 255;
assign img[15728] = 255;
assign img[15729] = 255;
assign img[15730] = 238;
assign img[15731] = 255;
assign img[15732] = 221;
assign img[15733] = 221;
assign img[15734] = 221;
assign img[15735] = 253;
assign img[15736] = 255;
assign img[15737] = 255;
assign img[15738] = 255;
assign img[15739] = 255;
assign img[15740] = 255;
assign img[15741] = 255;
assign img[15742] = 239;
assign img[15743] = 238;
assign img[15744] = 96;
assign img[15745] = 238;
assign img[15746] = 254;
assign img[15747] = 239;
assign img[15748] = 238;
assign img[15749] = 238;
assign img[15750] = 238;
assign img[15751] = 255;
assign img[15752] = 255;
assign img[15753] = 255;
assign img[15754] = 239;
assign img[15755] = 190;
assign img[15756] = 255;
assign img[15757] = 255;
assign img[15758] = 255;
assign img[15759] = 223;
assign img[15760] = 205;
assign img[15761] = 204;
assign img[15762] = 236;
assign img[15763] = 238;
assign img[15764] = 238;
assign img[15765] = 238;
assign img[15766] = 238;
assign img[15767] = 238;
assign img[15768] = 238;
assign img[15769] = 206;
assign img[15770] = 204;
assign img[15771] = 238;
assign img[15772] = 238;
assign img[15773] = 255;
assign img[15774] = 255;
assign img[15775] = 255;
assign img[15776] = 255;
assign img[15777] = 255;
assign img[15778] = 255;
assign img[15779] = 255;
assign img[15780] = 255;
assign img[15781] = 255;
assign img[15782] = 255;
assign img[15783] = 239;
assign img[15784] = 238;
assign img[15785] = 238;
assign img[15786] = 238;
assign img[15787] = 238;
assign img[15788] = 254;
assign img[15789] = 255;
assign img[15790] = 255;
assign img[15791] = 255;
assign img[15792] = 255;
assign img[15793] = 255;
assign img[15794] = 255;
assign img[15795] = 255;
assign img[15796] = 255;
assign img[15797] = 255;
assign img[15798] = 255;
assign img[15799] = 255;
assign img[15800] = 255;
assign img[15801] = 255;
assign img[15802] = 255;
assign img[15803] = 255;
assign img[15804] = 255;
assign img[15805] = 255;
assign img[15806] = 255;
assign img[15807] = 255;
assign img[15808] = 255;
assign img[15809] = 255;
assign img[15810] = 255;
assign img[15811] = 255;
assign img[15812] = 255;
assign img[15813] = 255;
assign img[15814] = 255;
assign img[15815] = 255;
assign img[15816] = 255;
assign img[15817] = 255;
assign img[15818] = 255;
assign img[15819] = 255;
assign img[15820] = 255;
assign img[15821] = 207;
assign img[15822] = 238;
assign img[15823] = 238;
assign img[15824] = 238;
assign img[15825] = 238;
assign img[15826] = 238;
assign img[15827] = 254;
assign img[15828] = 255;
assign img[15829] = 223;
assign img[15830] = 236;
assign img[15831] = 238;
assign img[15832] = 238;
assign img[15833] = 238;
assign img[15834] = 238;
assign img[15835] = 255;
assign img[15836] = 255;
assign img[15837] = 255;
assign img[15838] = 255;
assign img[15839] = 255;
assign img[15840] = 187;
assign img[15841] = 187;
assign img[15842] = 255;
assign img[15843] = 255;
assign img[15844] = 255;
assign img[15845] = 239;
assign img[15846] = 254;
assign img[15847] = 255;
assign img[15848] = 255;
assign img[15849] = 255;
assign img[15850] = 255;
assign img[15851] = 255;
assign img[15852] = 255;
assign img[15853] = 255;
assign img[15854] = 255;
assign img[15855] = 255;
assign img[15856] = 238;
assign img[15857] = 238;
assign img[15858] = 254;
assign img[15859] = 255;
assign img[15860] = 191;
assign img[15861] = 187;
assign img[15862] = 234;
assign img[15863] = 238;
assign img[15864] = 254;
assign img[15865] = 255;
assign img[15866] = 223;
assign img[15867] = 221;
assign img[15868] = 221;
assign img[15869] = 255;
assign img[15870] = 255;
assign img[15871] = 255;
assign img[15872] = 48;
assign img[15873] = 247;
assign img[15874] = 255;
assign img[15875] = 255;
assign img[15876] = 255;
assign img[15877] = 255;
assign img[15878] = 191;
assign img[15879] = 187;
assign img[15880] = 251;
assign img[15881] = 255;
assign img[15882] = 239;
assign img[15883] = 222;
assign img[15884] = 253;
assign img[15885] = 255;
assign img[15886] = 255;
assign img[15887] = 239;
assign img[15888] = 204;
assign img[15889] = 204;
assign img[15890] = 236;
assign img[15891] = 191;
assign img[15892] = 155;
assign img[15893] = 255;
assign img[15894] = 255;
assign img[15895] = 255;
assign img[15896] = 255;
assign img[15897] = 191;
assign img[15898] = 255;
assign img[15899] = 255;
assign img[15900] = 255;
assign img[15901] = 255;
assign img[15902] = 239;
assign img[15903] = 238;
assign img[15904] = 238;
assign img[15905] = 238;
assign img[15906] = 238;
assign img[15907] = 238;
assign img[15908] = 238;
assign img[15909] = 254;
assign img[15910] = 254;
assign img[15911] = 255;
assign img[15912] = 238;
assign img[15913] = 238;
assign img[15914] = 238;
assign img[15915] = 238;
assign img[15916] = 238;
assign img[15917] = 238;
assign img[15918] = 238;
assign img[15919] = 238;
assign img[15920] = 254;
assign img[15921] = 255;
assign img[15922] = 255;
assign img[15923] = 255;
assign img[15924] = 255;
assign img[15925] = 255;
assign img[15926] = 255;
assign img[15927] = 255;
assign img[15928] = 255;
assign img[15929] = 255;
assign img[15930] = 255;
assign img[15931] = 255;
assign img[15932] = 255;
assign img[15933] = 255;
assign img[15934] = 255;
assign img[15935] = 255;
assign img[15936] = 255;
assign img[15937] = 255;
assign img[15938] = 255;
assign img[15939] = 255;
assign img[15940] = 255;
assign img[15941] = 255;
assign img[15942] = 255;
assign img[15943] = 239;
assign img[15944] = 238;
assign img[15945] = 238;
assign img[15946] = 254;
assign img[15947] = 255;
assign img[15948] = 255;
assign img[15949] = 255;
assign img[15950] = 255;
assign img[15951] = 255;
assign img[15952] = 255;
assign img[15953] = 255;
assign img[15954] = 255;
assign img[15955] = 255;
assign img[15956] = 255;
assign img[15957] = 255;
assign img[15958] = 255;
assign img[15959] = 255;
assign img[15960] = 239;
assign img[15961] = 238;
assign img[15962] = 238;
assign img[15963] = 238;
assign img[15964] = 238;
assign img[15965] = 238;
assign img[15966] = 238;
assign img[15967] = 191;
assign img[15968] = 239;
assign img[15969] = 238;
assign img[15970] = 238;
assign img[15971] = 238;
assign img[15972] = 238;
assign img[15973] = 238;
assign img[15974] = 190;
assign img[15975] = 187;
assign img[15976] = 251;
assign img[15977] = 255;
assign img[15978] = 255;
assign img[15979] = 255;
assign img[15980] = 221;
assign img[15981] = 255;
assign img[15982] = 255;
assign img[15983] = 255;
assign img[15984] = 221;
assign img[15985] = 221;
assign img[15986] = 221;
assign img[15987] = 255;
assign img[15988] = 221;
assign img[15989] = 221;
assign img[15990] = 253;
assign img[15991] = 255;
assign img[15992] = 255;
assign img[15993] = 191;
assign img[15994] = 234;
assign img[15995] = 174;
assign img[15996] = 170;
assign img[15997] = 238;
assign img[15998] = 238;
assign img[15999] = 238;
assign img[16000] = 96;
assign img[16001] = 255;
assign img[16002] = 255;
assign img[16003] = 223;
assign img[16004] = 204;
assign img[16005] = 204;
assign img[16006] = 204;
assign img[16007] = 236;
assign img[16008] = 238;
assign img[16009] = 239;
assign img[16010] = 238;
assign img[16011] = 206;
assign img[16012] = 204;
assign img[16013] = 220;
assign img[16014] = 157;
assign img[16015] = 187;
assign img[16016] = 234;
assign img[16017] = 255;
assign img[16018] = 255;
assign img[16019] = 255;
assign img[16020] = 238;
assign img[16021] = 238;
assign img[16022] = 238;
assign img[16023] = 255;
assign img[16024] = 254;
assign img[16025] = 255;
assign img[16026] = 255;
assign img[16027] = 255;
assign img[16028] = 255;
assign img[16029] = 255;
assign img[16030] = 255;
assign img[16031] = 255;
assign img[16032] = 238;
assign img[16033] = 254;
assign img[16034] = 255;
assign img[16035] = 255;
assign img[16036] = 255;
assign img[16037] = 255;
assign img[16038] = 255;
assign img[16039] = 255;
assign img[16040] = 238;
assign img[16041] = 238;
assign img[16042] = 255;
assign img[16043] = 255;
assign img[16044] = 239;
assign img[16045] = 238;
assign img[16046] = 238;
assign img[16047] = 238;
assign img[16048] = 238;
assign img[16049] = 255;
assign img[16050] = 255;
assign img[16051] = 255;
assign img[16052] = 255;
assign img[16053] = 255;
assign img[16054] = 255;
assign img[16055] = 255;
assign img[16056] = 255;
assign img[16057] = 255;
assign img[16058] = 239;
assign img[16059] = 238;
assign img[16060] = 238;
assign img[16061] = 255;
assign img[16062] = 255;
assign img[16063] = 255;
assign img[16064] = 255;
assign img[16065] = 255;
assign img[16066] = 255;
assign img[16067] = 255;
assign img[16068] = 255;
assign img[16069] = 255;
assign img[16070] = 238;
assign img[16071] = 254;
assign img[16072] = 255;
assign img[16073] = 255;
assign img[16074] = 255;
assign img[16075] = 255;
assign img[16076] = 255;
assign img[16077] = 255;
assign img[16078] = 255;
assign img[16079] = 255;
assign img[16080] = 255;
assign img[16081] = 255;
assign img[16082] = 255;
assign img[16083] = 255;
assign img[16084] = 238;
assign img[16085] = 238;
assign img[16086] = 238;
assign img[16087] = 255;
assign img[16088] = 238;
assign img[16089] = 238;
assign img[16090] = 238;
assign img[16091] = 238;
assign img[16092] = 254;
assign img[16093] = 255;
assign img[16094] = 255;
assign img[16095] = 255;
assign img[16096] = 238;
assign img[16097] = 238;
assign img[16098] = 238;
assign img[16099] = 238;
assign img[16100] = 238;
assign img[16101] = 238;
assign img[16102] = 238;
assign img[16103] = 238;
assign img[16104] = 238;
assign img[16105] = 255;
assign img[16106] = 255;
assign img[16107] = 255;
assign img[16108] = 239;
assign img[16109] = 255;
assign img[16110] = 255;
assign img[16111] = 255;
assign img[16112] = 255;
assign img[16113] = 255;
assign img[16114] = 187;
assign img[16115] = 223;
assign img[16116] = 221;
assign img[16117] = 221;
assign img[16118] = 204;
assign img[16119] = 238;
assign img[16120] = 238;
assign img[16121] = 223;
assign img[16122] = 221;
assign img[16123] = 205;
assign img[16124] = 220;
assign img[16125] = 253;
assign img[16126] = 255;
assign img[16127] = 255;
assign img[16128] = 64;
assign img[16129] = 254;
assign img[16130] = 255;
assign img[16131] = 223;
assign img[16132] = 221;
assign img[16133] = 255;
assign img[16134] = 223;
assign img[16135] = 253;
assign img[16136] = 255;
assign img[16137] = 255;
assign img[16138] = 255;
assign img[16139] = 255;
assign img[16140] = 204;
assign img[16141] = 236;
assign img[16142] = 238;
assign img[16143] = 238;
assign img[16144] = 204;
assign img[16145] = 236;
assign img[16146] = 238;
assign img[16147] = 238;
assign img[16148] = 220;
assign img[16149] = 253;
assign img[16150] = 255;
assign img[16151] = 255;
assign img[16152] = 255;
assign img[16153] = 255;
assign img[16154] = 223;
assign img[16155] = 204;
assign img[16156] = 252;
assign img[16157] = 255;
assign img[16158] = 255;
assign img[16159] = 255;
assign img[16160] = 255;
assign img[16161] = 255;
assign img[16162] = 255;
assign img[16163] = 255;
assign img[16164] = 255;
assign img[16165] = 255;
assign img[16166] = 255;
assign img[16167] = 255;
assign img[16168] = 255;
assign img[16169] = 255;
assign img[16170] = 239;
assign img[16171] = 238;
assign img[16172] = 254;
assign img[16173] = 239;
assign img[16174] = 238;
assign img[16175] = 255;
assign img[16176] = 255;
assign img[16177] = 255;
assign img[16178] = 255;
assign img[16179] = 255;
assign img[16180] = 255;
assign img[16181] = 255;
assign img[16182] = 255;
assign img[16183] = 255;
assign img[16184] = 255;
assign img[16185] = 255;
assign img[16186] = 255;
assign img[16187] = 255;
assign img[16188] = 255;
assign img[16189] = 207;
assign img[16190] = 238;
assign img[16191] = 255;
assign img[16192] = 255;
assign img[16193] = 255;
assign img[16194] = 223;
assign img[16195] = 255;
assign img[16196] = 255;
assign img[16197] = 255;
assign img[16198] = 255;
assign img[16199] = 255;
assign img[16200] = 255;
assign img[16201] = 255;
assign img[16202] = 255;
assign img[16203] = 255;
assign img[16204] = 223;
assign img[16205] = 255;
assign img[16206] = 255;
assign img[16207] = 255;
assign img[16208] = 255;
assign img[16209] = 255;
assign img[16210] = 255;
assign img[16211] = 239;
assign img[16212] = 238;
assign img[16213] = 239;
assign img[16214] = 238;
assign img[16215] = 238;
assign img[16216] = 254;
assign img[16217] = 255;
assign img[16218] = 255;
assign img[16219] = 255;
assign img[16220] = 255;
assign img[16221] = 255;
assign img[16222] = 255;
assign img[16223] = 239;
assign img[16224] = 220;
assign img[16225] = 253;
assign img[16226] = 255;
assign img[16227] = 255;
assign img[16228] = 223;
assign img[16229] = 221;
assign img[16230] = 221;
assign img[16231] = 221;
assign img[16232] = 252;
assign img[16233] = 255;
assign img[16234] = 255;
assign img[16235] = 255;
assign img[16236] = 255;
assign img[16237] = 237;
assign img[16238] = 238;
assign img[16239] = 206;
assign img[16240] = 204;
assign img[16241] = 220;
assign img[16242] = 253;
assign img[16243] = 223;
assign img[16244] = 205;
assign img[16245] = 204;
assign img[16246] = 236;
assign img[16247] = 238;
assign img[16248] = 238;
assign img[16249] = 238;
assign img[16250] = 238;
assign img[16251] = 255;
assign img[16252] = 255;
assign img[16253] = 255;
assign img[16254] = 255;
assign img[16255] = 239;
assign img[16256] = 96;
assign img[16257] = 70;
assign img[16258] = 100;
assign img[16259] = 238;
assign img[16260] = 238;
assign img[16261] = 238;
assign img[16262] = 238;
assign img[16263] = 222;
assign img[16264] = 238;
assign img[16265] = 255;
assign img[16266] = 206;
assign img[16267] = 206;
assign img[16268] = 254;
assign img[16269] = 255;
assign img[16270] = 221;
assign img[16271] = 205;
assign img[16272] = 204;
assign img[16273] = 204;
assign img[16274] = 252;
assign img[16275] = 239;
assign img[16276] = 138;
assign img[16277] = 200;
assign img[16278] = 200;
assign img[16279] = 254;
assign img[16280] = 255;
assign img[16281] = 255;
assign img[16282] = 255;
assign img[16283] = 255;
assign img[16284] = 255;
assign img[16285] = 255;
assign img[16286] = 239;
assign img[16287] = 238;
assign img[16288] = 204;
assign img[16289] = 253;
assign img[16290] = 255;
assign img[16291] = 255;
assign img[16292] = 239;
assign img[16293] = 238;
assign img[16294] = 255;
assign img[16295] = 255;
assign img[16296] = 238;
assign img[16297] = 238;
assign img[16298] = 255;
assign img[16299] = 255;
assign img[16300] = 255;
assign img[16301] = 255;
assign img[16302] = 238;
assign img[16303] = 238;
assign img[16304] = 254;
assign img[16305] = 255;
assign img[16306] = 255;
assign img[16307] = 239;
assign img[16308] = 238;
assign img[16309] = 255;
assign img[16310] = 238;
assign img[16311] = 255;
assign img[16312] = 255;
assign img[16313] = 255;
assign img[16314] = 255;
assign img[16315] = 255;
assign img[16316] = 255;
assign img[16317] = 239;
assign img[16318] = 238;
assign img[16319] = 255;
assign img[16320] = 255;
assign img[16321] = 255;
assign img[16322] = 255;
assign img[16323] = 255;
assign img[16324] = 255;
assign img[16325] = 255;
assign img[16326] = 255;
assign img[16327] = 255;
assign img[16328] = 239;
assign img[16329] = 238;
assign img[16330] = 238;
assign img[16331] = 223;
assign img[16332] = 221;
assign img[16333] = 253;
assign img[16334] = 255;
assign img[16335] = 255;
assign img[16336] = 255;
assign img[16337] = 255;
assign img[16338] = 239;
assign img[16339] = 238;
assign img[16340] = 238;
assign img[16341] = 238;
assign img[16342] = 238;
assign img[16343] = 238;
assign img[16344] = 238;
assign img[16345] = 238;
assign img[16346] = 238;
assign img[16347] = 238;
assign img[16348] = 238;
assign img[16349] = 174;
assign img[16350] = 186;
assign img[16351] = 239;
assign img[16352] = 204;
assign img[16353] = 204;
assign img[16354] = 252;
assign img[16355] = 255;
assign img[16356] = 255;
assign img[16357] = 255;
assign img[16358] = 174;
assign img[16359] = 254;
assign img[16360] = 255;
assign img[16361] = 239;
assign img[16362] = 238;
assign img[16363] = 255;
assign img[16364] = 239;
assign img[16365] = 255;
assign img[16366] = 223;
assign img[16367] = 221;
assign img[16368] = 221;
assign img[16369] = 221;
assign img[16370] = 221;
assign img[16371] = 221;
assign img[16372] = 255;
assign img[16373] = 255;
assign img[16374] = 255;
assign img[16375] = 255;
assign img[16376] = 223;
assign img[16377] = 221;
assign img[16378] = 253;
assign img[16379] = 239;
assign img[16380] = 238;
assign img[16381] = 238;
assign img[16382] = 255;
assign img[16383] = 255;
end

endmodule
