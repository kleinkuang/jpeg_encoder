// File:    jpeg_encoder_tb.sv
// Author:  Lei Kuang
// Date:    15th July 2020
// @ Imperial College London

module jpeg_encoder_tb;

logic        clk;
logic        nrst;

logic [7:0]  din;
logic        din_valid;
logic [31:0] dout;
logic        dout_valid;

jpeg_encoder dut(.*);

initial begin
    clk = '0;
    forever #5ns clk = ~clk;
end

logic [7:0]  seq [0:16383];
logic [13:0] cnt;

logic [7:0] cnt_t = '0;

always_ff @ (posedge clk)
    //cnt_t <= cnt_t + 1;
    cnt_t <= '1;
    
assign din_valid = cnt_t=='1;

initial begin
    nrst      = '0;
    cnt       = '0;
    //din_valid = '0;

    @(posedge clk)
        nrst <= '1;
    
    forever begin
        @(posedge clk) begin
            //din_valid <= ~din_valid;
            
            if(din_valid)
                cnt <= cnt + 1;
        end
    end
end

always_ff @ (negedge clk)
    if(dout_valid)
        $write("%8X\n", dout);

assign din = seq[cnt];

assign seq = '{

  45, -19,   3,  -1,   1, -19, -13,   1,
  -3,   3,   0,   2,  -3,   2,  -7,  -3,
   0,   0,   0,   1,   2,  -2,   0,  -1,
   0,   0,   0,  -1,  -1,   0,   0,   1,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   4,   0,  -1,   1,  -1,   1,   0,
   0,   1,   0,   1,  -1,  -1,  -2,   0,
   0,   1,  -2,  -1,  -1,  -1,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,  -8,  -1,   1,  -1,  -1,  -3,   0,
   0,  -3,   2,   0,   2,  -1,  -1,   0,
  -1,  -1,   1,   0,  -1,   0,   1,  -1,
  -1,  -1,   0,   1,   0,   0,   0,   0,
   0,   1,   0,   1,   0,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   1,   1,   1,   0,   0,   4,   1,
  -1,  -3,   0,   1,  -1,   0,   0,   0,
   0,  -1,   0,   0,   0,   0,  -2,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,  -1,  -2,   0,   0,  -3,  -2,   3,
  -1,  -1,  -1,  -1,   1,   1,  -1,   0,
   1,   1,  -1,   0,   1,   0,   0,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   1,   0,   1,   0,   2,   0,   2,
  -2,   0,  -3,   1,  -1,   0,   0,   0,
   1,  -1,   0,   1,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,   0,   1,  -1,   2,   1,   0,  -1,
   1,   0,  -1,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   1,  -2,   1,  -1,   2,   0,   2,
   1,   3,   1,   1,  -1,   1,   1,  -1,
   0,  -2,  -1,   0,  -1,   0,   0,  -1,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   3,  -3,   3,   1,   2,  -1,   1,
   0,   3,   2,   0,  -1,  -1,   1,   0,
   1,   1,   0,   0,  -2,  -1,   0,   0,
   1,   0,   0,   0,   0,   0,   0,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,  -2,   0,   0,   0,   1,   0,   0,
   0,   0,  -1,   0,  -2,   0,   0,   0,
   0,  -1,  -1,  -1,  -1,   0,   0,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   1,   1,  -1,   0,   0,   0,   1,
   1,  -1,   0,  -1,   1,   1,   0,   0,
   1,   0,   0,   0,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,  -2,   1,  -2,   5,  -3,   0,   1,
   0,   0,   0,   1,  -1,   2,  -1,   0,
   0,   0,  -1,   1,   1,   1,   0,   0,
   1,  -1,   0,   0,   0,   0,   0,   0,
   0,  -1,   1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -3,  -3,  -2,   3,  -7,  -3,   1,
  -3,  -1,  -1,   0,   0,   0,   0,  -1,
   1,  -2,   2,  -1,   0,  -1,   0,   0,
   0,   0,   0,   1,   0,   0,  -1,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   0,  -2,   3,  -1,   1,   0,   0,
  -1,   0,  -1,   1,  -1,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,  -1,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,  -8,   1,   0,   1,  -3,  -3,   0,
   1,   0,   0,   1,   3,   0,  -1,   1,
  -1,   1,   0,   0,   1,   0,  -1,   0,
  -1,   0,   0,   0,   0,   0,   0,  -1,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,  -3,  -3,  -2,  -3,   3,   1,   0,
  -2,   1,   1,   0,  -2,   1,  -1,   1,
   1,   1,  -1,   2,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  43, -16,  -5,   0,   2, -16, -13,   0,
  -2,   2,   1,  -1,  -1,   0,  -5,  -2,
   0,   0,   1,   0,  -1,  -1,   0,   1,
   0,   1,   0,  -1,   0,   0,   0,   0,
   0,   1,   1,  -1,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  51,   3,  -1,  -4,  -3,   7,   2,   1,
   1,   2,  -3,  -2,   3,   0,  -1,   0,
   1,   1,   0,  -1,  -3,  -1,  -1,   1,
   1,   0,  -1,   0,   0,   0,   0,   0,
   1,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  53,  -5,   2,   2,   2,   2,  -1,   2,
   4,   2,   3,   0,   2,   2,   0,   0,
  -1,  -1,  -1,  -2,  -1,   1,   1,  -2,
  -1,  -1,   0,   1,   0,   0,   0,   0,
   0,   1,  -1,   0,   0,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,  -3,  -2,  -2,  -3,   0,   6,  -2,
   2,   2,  -2,  -2,   0,   1,   1,   1,
   1,   0,   1,  -1,   0,   0,   0,   0,
   0,   0,   1,   0,  -1,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  53,  -7,   1,   5,  -2,  -5,  -4,   0,
   3,  -5,  -2,  -1,   0,   0,   0,   0,
   0,   0,   0,  -2,   0,   0,  -1,  -1,
  -1,  -1,   0,  -1,   0,   0,   0,   0,
   0,  -1,   0,   1,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   3,   0,  -2,   5,   0,   1,  -2,
  -1,   1,   0,   0,   2,   0,  -1,   0,
   0,  -1,   0,   0,   1,   0,   0,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,  -1,  -4,  -1,  -1,   2,   0,   2,
   1,   0,   1,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   2,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,  -1,  -1,   0,  -1,   2,   0,  -1,
   1,   0,   0,   0,   0,   0,   1,   0,
   1,   0,   0,   0,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,   4,   2,   2,  -1,  -1,   0,   0,
  -2,  -2,  -1,   1,   0,   0,   1,   0,
  -1,   1,   0,   1,   1,   0,  -1,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,  -1,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,  -1,  -1,   1,   0,   1,  -1,   1,
   2,   1,  -1,   0,   0,   1,  -1,   0,
   0,   1,  -1,  -1,   1,   0,   0,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   3,   2,  -1,   1,   3,  -1,  -1,
   0,   1,  -1,   0,   0,   1,   0,   0,
   0,  -1,   0,   0,  -1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,   3,   0,   1,   1,  -3,   1,  -1,
  -1,   2,  -2,   1,  -1,   0,  -2,   0,
   0,   1,   1,   1,   1,   1,   0,  -1,
   0,   0,   0,   0,   1,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -3,  -1,  -1,   2,  -8,  -4,   0,
  -2,   2,  -1,   5,  -2,   0,   1,  -1,
   0,   0,   1,   1,   1,   1,   0,  -1,
   1,   0,   0,   1,   0,   0,   0,   0,
   0,   1,   1,   0,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   1,   0,   0,   1,   1,   1,  -2,
   0,   0,   1,  -2,   1,   0,  -1,   0,
   0,  -1,   1,   0,  -2,   0,   0,  -1,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,  -2,   3,  -1,   2,   0,   0,   0,
   1,   5,  -2,   2,   2,   0,   0,   0,
   0,   0,   0,   0,  -1,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,  -3,  -2,   1,   2,   2,   1,  -2,
   1,  -1,   1,   0,   0,  -1,   1,   0,
   1,   0,   1,   0,  -1,  -1,  -1,   0,
   0,   0,   0,   1,   0,   0,   0,   0,
   0,   0,  -1,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  43, -23,   1,   1,   2, -19, -12,   1,
   3,   2,   1,   0,  -1,   1,  -5,  -2,
   1,  -2,   0,  -1,  -1,   1,  -3,  -1,
   0,  -1,   0,  -1,  -1,   0,  -1,   0,
   1,   0,   0,   0,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,   6,  -2,   1,   1,   1,   0,  -2,
   2,  -1,  -1,   0,  -2,   0,  -1,   0,
   0,   1,   2,   0,   2,   1,  -1,   0,
  -1,   0,   0,   0,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   1,   0,
   0,   0,   0,   0,   0,   0,  -1,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  51,  -3,   2,   6,  -3,   2,  -3,  -4,
  -1,  -2,  -5,   0,   0,  -2,  -2,   0,
   0,   1,   2,   1,   3,   0,   0,   1,
   0,   0,   0,   1,   0,   0,   1,   0,
   0,   0,  -1,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -3,   2,   2,   3,   0,   5,   0,
   1,  -1,   2,  -1,   1,  -1,   1,   0,
  -1,  -1,   0,   1,   0,   0,   0,   0,
   1,  -1,   0,  -1,  -1,   0,   0,   0,
  -1,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,  -4,  -2,  -2,  -1,  -9,  -4,   0,
  -3,   2,   0,  -2,  -4,  -1,  -3,  -1,
   0,  -1,   0,   0,  -1,   0,   0,   0,
  -1,  -1,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,  -2,  -4,  -3,  -2,   4,   1,   2,
   0,  -2,  -1,   0,   3,   2,   1,   0,
  -1,   1,   1,   1,   0,   0,   0,   1,
   0,   0,   0,  -1,  -1,   0,   0,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  62,   0,   0,  -1,  -2,   0,   0,   1,
   0,   0,  -1,  -1,  -1,   0,   0,   0,
   0,   1,   0,   0,  -1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,  -2,   2,  -1,   0,   1,   0,   1,
   1,   0,   0,   0,   0,   1,   1,   0,
   0,  -1,   0,   0,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   3,   2,   0,  -1,  -1,   1,   0,
   2,   0,   1,  -1,  -1,   0,   0,   0,
   0,   0,   1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,  -2,   2,  -2,   1,   0,  -1,  -1,
  -1,  -1,   0,   1,  -1,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,   2,   1,  -1,   3,   3,   0,   2,
   2,   0,  -2,   0,  -1,  -3,   1,   0,
   0,  -1,  -1,   0,   1,   0,   0,   1,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,  -1,   0,  -1,   1,  -5,   2,   2,
  -2,   0,   0,   2,  -2,   1,  -1,   0,
   0,   0,  -1,  -2,   2,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
  -1,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,  -1,  -4,  -1,  -4, -10,  -3,  -3,
  -2,   4,   1,  -1,  -2,  -1,   1,   0,
  -1,  -1,   2,   0,   0,  -1,   1,   1,
   0,   0,   1,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,   1,   2,   0,  -1,   4,   1,  -1,
   1,  -1,  -3,   1,   2,   0,  -1,   1,
   0,  -1,   0,   0,   0,  -1,   0,   2,
   2,   0,   0,   0,   0,   0,   0,   0,
  -1,  -1,   0,   0,   0,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  47,  -8,   0,   1,  -1,   4,  -1,   1,
   1,  -5,   5,   0,  -2,   0,   0,   0,
   0,  -1,   2,   4,   4,   0,   1,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,  -1,  -1,   1,   1,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,  -2,  -2,  -1,  -2,   1,   2,   1,
  -3,  -2,  -3,   0,   2,   3,   1,   0,
   1,   2,   0,  -2,   0,   0,   0,   0,
   1,   0,   0,   1,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  43, -23,   0,   0,  -6, -24, -14,  -3,
   3,   1,  -4,  -3,   2,   0,  -6,  -3,
   0,   0,  -2,  -3,  -1,   0,   0,  -1,
   0,   0,   0,  -1,   0,   0,   0,   0,
  -1,   0,   0,   0,  -1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,   0,  -3,  -1,   0,   2,   0,   2,
   0,   2,  -1,   0,  -1,   0,  -1,   0,
   0,   0,   1,   0,  -2,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,  -2,   2,   0,  -2,   2,  -2,  -1,
   2,  -1,   2,   0,  -1,   0,  -2,   0,
   0,   0,   3,   1,   0,   0,   0,   0,
   0,   0,   0,   1,   0,   0,  -1,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  53,  -2,  -1,  -4,  -2,   1,   7,   2,
   1,  -2,  -1,  -1,  -1,   1,   1,   0,
   1,   1,   0,  -1,  -2,  -1,  -1,   1,
   2,   0,   0,   0,   0,   0,   0,   0,
   0,   1,   0,   0,   0,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   1,   0,

  59,  -3,   1,   0,   3,  -6,  -2,   1,
  -2,   1,   1,  -3,   1,   2,  -2,   0,
   1,   0,   0,   1,  -1,  -1,   0,   1,
  -1,   1,   0,   0,   0,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,   0,  -2,  -2,   1,   6,   2,  -2,
   3,   2,   0,   0,   1,   0,  -1,   0,
   1,  -1,   0,   0,   1,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,  -1,  -3,  -1,  -1,   1,   0,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,   1,  -1,  -1,   0,   1,  -1,   1,
   0,   1,   1,   0,  -1,   0,   2,   0,
   1,   0,   0,   0,   1,   0,   1,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,   2,   0,   0,   0,   0,   0,   1,
  -1,  -1,   0,   1,   1,   0,   1,   0,
   0,   1,   0,   0,   0,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,   1,   1,   1,  -1,   1,  -1,  -1,
   0,  -1,   1,   0,   0,   0,   0,   0,
   0,   0,   1,   0,   0,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   0,   0,  -2,  -2,   2,  -2,  -2,
   0,   1,   0,   0,  -1,   0,   0,   0,
  -1,  -1,   0,   0,  -1,   1,   1,  -1,
  -1,   0,   0,   0,   0,   0,   0,   0,
   1,   1,   0,   0,   0,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,  -2,   1,   1,   1,  -2,   0,   0,
  -1,   2,   0,   1,   0,  -1,   0,   0,
   0,   0,   0,   0,  -2,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,   1,   0,   1,   3,  -8,  -2,   3,
  -2,  -4,  -1,   0,   1,   0,   1,   0,
   1,   0,  -2,   4,   0,   1,   0,   0,
  -1,   0,   0,   1,   0,   0,   0,   0,
   0,   0,   0,  -1,   0,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   3,  -1,  -2,   2,   0,  -1,   1,
   1,  -1,  -1,   0,   2,   0,  -1,   1,
  -1,   0,   0,   0,   1,  -1,   0,   1,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,  -3,  -3,  -2,   2,   1,  -2,   2,
   2,   0,  -1,   1,   1,  -1,  -1,   0,
  -1,   0,   0,   2,   0,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,  -3,  -3,  -2,  -1,   6,   3,   1,
  -2,  -1,  -2,  -2,   3,   2,   0,   0,
   1,   2,  -1,  -1,   2,   1,   0,   0,
   1,   0,   0,   0,   0,   0,  -1,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  41, -14,   1,  -6,   0, -18, -14,   0,
   4,   3,  -2,  -2,   0,   2,  -5,  -2,
  -1,  -1,  -3,   2,  -1,  -1,   0,  -1,
   2,   0,   0,   0,  -1,   0,   0,  -1,
   0,  -1,   1,  -1,   0,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,   5,  -3,  -1,   1,   2,   0,   0,
  -1,  -1,   2,  -1,   0,   0,  -2,   0,
   0,  -1,   2,  -1,   1,   1,  -1,   0,
   0,   1,   0,   0,   0,   0,  -1,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   2,   2,   1,   2,   5,  -2,  -3,
   1,  -1,   1,  -1,   1,   1,  -2,   0,
   2,   0,   0,   1,   0,  -1,   0,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   0,   0,  -2,   1,  -1,   3,  -2,
   4,  -1,  -2,  -2,  -1,   1,  -1,   0,
  -1,   2,  -1,   0,   1,   0,   0,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   1,   0,   0,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,  -5,  -1,   1,  -1,  -4,  -2,   0,
   1,  -1,   0,  -1,   0,   0,  -1,   0,
   1,   1,   0,   2,  -1,   0,   0,   0,
  -1,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,  -1,  -1,   1,   1,   1,   0,   0,
   1,  -1,   1,  -1,   1,   0,   0,   0,
   0,   0,   1,   0,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  63,   0,   1,   0,   0,   1,   0,  -1,
   0,   1,  -1,   0,   0,   0,   0,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   3,   2,   1,  -2,   5,  -2,   1,
  -2,   1,  -1,   0,   0,   2,   2,   0,
  -1,   2,   0,   1,   1,   0,   0,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   1,   0,   1,   1,   3,   2,   0,
   2,   0,   0,  -1,  -2,  -1,   1,   0,
   0,  -1,   0,   0,   2,   0,   0,   0,
   1,   0,   0,  -1,   0,   0,   0,  -1,
   1,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,  -1,   0,   0,   2,   0,  -1,   2,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,  -1,   1,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   1,   1,  -1,   0,   1,  -1,  -2,
   1,   1,   1,   0,  -2,   0,   0,   0,
   0,   0,   0,  -1,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   3,   1,   1,  -1,  -8,   2,  -1,
   1,   1,   1,   0,  -1,   0,  -3,   0,
   0,   0,   1,   0,   1,   0,   0,   1,
   1,  -1,   0,  -1,   0,   0,   0,   1,
   0,   1,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -3,   1,  -2,  -1, -10,  -2,   1,
  -3,   1,  -2,  -1,  -2,  -2,   0,   0,
  -1,   0,   1,   0,   2,   0,   1,  -1,
   0,   0,   0,   1,   0,   0,   0,  -1,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   2,  -2,   0,   1,   0,   0,   0,
   0,  -1,   1,  -1,  -1,   0,  -1,   0,
  -1,   1,   1,  -1,   1,   0,  -1,   1,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,  -2,  -7,  -2,  -4,   4,  -1,   0,
  -2,   0,   1,   1,   0,   0,  -1,   0,
   0,   0,   1,   1,   1,   1,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,  -1,   0,   1,   0,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,  -2,  -3,   1,  -2,   2,   2,   1,
   1,   1,   1,   0,  -2,   0,   1,   0,
   0,  -1,  -2,   0,  -1,   0,  -1,  -1,
   0,   0,   0,   0,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   1,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  44, -16,  -2,  -1,   0, -18, -11,   3,
  -2,  -1,   0,   0,   2,  -1,  -7,  -2,
   0,   0,   0,   1,  -1,   2,   2,   0,
   0,   0,   0,  -1,  -1,   0,   0,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,  -1,   0,   0,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  51,   8,   1,  -1,  -1,   3,   1,   0,
   2,   0,  -1,   0,  -4,  -1,  -2,   0,
   0,   2,   1,   1,   0,   0,  -2,   0,
  -1,   0,   0,   0,   0,   0,   0,   1,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  53,  -7,  -3,   0,  -4,   0,  -3,   0,
  -2,   0,   0,  -1,  -1,  -1,  -2,   0,
  -1,  -1,  -3,  -1,  -2,   0,  -1,   0,
   0,   0,   0,   1,   0,   0,   0,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -1,   3,   1,   3,  -4,   7,   1,
   0,  -4,  -1,  -1,   0,   0,   0,   1,
  -1,   0,  -1,  -1,   0,   0,   0,   0,
   2,   0,   0,  -1,   0,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,  -1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,  -3,   0,   0,   1,  -4,  -3,   2,
  -1,   0,   3,  -2,   0,  -1,  -2,   0,
   0,   0,  -2,   0,  -1,   0,  -1,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,   2,   3,  -3,   1,   0,  -1,  -2,
   1,   2,   0,  -1,   1,   1,   1,   0,
   0,  -1,  -1,   0,   1,   1,   0,   0,
   0,   1,  -1,   0,   0,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,  -1,   0,   2,   1,   1,  -1,   1,
   1,   0,   0,  -1,   0,   0,  -1,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,  -1,   2,  -1,   0,   1,   0,   0,
   1,   1,   0,   1,   0,   1,   2,  -1,
  -1,   1,   1,   0,  -1,  -1,   1,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,   0,  -3,  -2,   1,   1,   2,   0,
  -1,   0,  -2,   1,   0,   0,   1,   0,
   0,   1,  -1,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,  -1,   1,   0,  -1,  -1,  -1,  -1,
  -1,   0,  -1,  -1,   1,   0,   0,   0,
   0,   0,  -1,   1,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,   1,  -1,  -2,  -3,   3,   0,  -3,
  -1,   0,   1,  -2,   1,   1,   0,   0,
   0,  -1,  -1,   1,   2,   0,   0,   0,
   1,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,  -1,   1,  -1,   1,  -4,   1,   0,
   0,   2,   0,   2,  -1,   1,  -2,   0,
   0,   0,  -1,   0,   1,   0,   1,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,  -4,   2,  -1,  -1,  -8,  -3,   0,
  -1,  -1,   1,  -3,  -1,   0,   1,   0,
   0,   0,  -2,   2,   0,  -1,  -1,   1,
   0,   0,   0,   1,   0,   0,   0,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,   4,   1,   1,   1,   4,  -2,  -1,
  -2,   0,  -1,   0,  -1,  -1,  -1,   1,
   0,   1,  -1,   2,  -1,   1,   0,   0,
   1,   0,   0,   0,   0,   0,  -1,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  51,  -5,   0,   2,   1,   1,  -2,   0,
  -3,  -5,  -1,  -1,  -3,   0,   1,   0,
   0,   0,   2,  -1,   1,   0,   1,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,  -1,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  53,  -3,  -3,  -3,  -3,  10,   4,   3,
   0,   6,   1,   1,   1,   2,   0,  -1,
   0,   1,  -1,   0,  -1,  -1,   0,   0,
  -1,   0,  -1,   0,   0,   0,  -1,  -1,
   0,   1,  -1,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  44, -20,   0,   0,  -2, -17, -12,   0,
  -1,  -2,   0,   0,   2,   1,  -5,  -2,
   0,   0,  -1,   0,   1,   1,   0,   0,
   1,  -1,   0,   0,  -1,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  53,   4,   0,  -2,  -2,   5,  -1,   4,
   1,  -5,  -1,  -1,   2,   1,  -2,   0,
  -1,   0,   2,  -1,  -1,   0,   0,   2,
   0,   0,   0,   0,  -1,   0,   0,  -1,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  53,   0,  -2,  -4,  -2,   3,  -2,  -2,
   1,   0,  -1,   0,   4,   1,  -2,   0,
   0,   0,   2,  -1,  -2,   0,   0,   0,
   0,  -1,   0,   1,  -1,   0,   0,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -3,  -3,  -1,   1,   0,   5,  -1,
   2,   1,  -2,   4,  -1,   0,   1,   0,
   0,   1,  -1,   0,  -1,   0,   0,   0,
  -1,   0,   0,  -1,  -1,   0,   0,  -1,
   1,   0,   0,   0,   0,  -1,   0,   0,
   0,  -1,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -7,  -4,  -2,  -6, -10,  -5,  -2,
  -1,   0,   2,   0,  -1,   0,  -2,  -1,
  -1,   0,   1,   0,   0,   1,   0,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,  -2,   0,   1,   0,   0,   0,   0,
  -2,   1,  -1,   1,  -1,   0,   1,   0,
  -1,   0,   0,   1,   0,   0,  -1,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,  -1,  -1,   0,   0,   2,   0,   0,
  -1,   2,  -1,   1,   0,   0,   0,   0,
   1,   1,   0,  -1,   0,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   0,  -2,  -1,  -2,   1,  -1,   1,
   0,   0,   2,  -1,   2,   2,   1,   0,
   0,  -1,   0,   0,   1,   1,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   1,  -1,   2,   0,   0,   0,   0,
   2,   1,   0,   0,   0,  -1,   2,   0,
   0,   0,   0,  -1,   1,   1,  -1,   0,
   0,  -1,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,   0,  -1,  -1,   1,  -1,  -1,   1,
   1,   1,   0,   1,  -1,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   0,   2,   0,   1,   0,  -1,  -2,
   0,   2,   0,   1,   0,  -1,   1,   0,
  -1,   1,   1,   0,   0,   1,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   3,  -1,   3,   1,  -4,   1,   1,
   0,   0,  -1,  -1,   1,   0,  -2,   1,
   0,   0,   0,   0,   0,   1,   0,   0,
  -1,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,  -2,  -1,  -2,  -3,  -3,  -1,  -3,
  -3,   0,   0,  -1,  -1,  -1,   0,   0,
   0,   0,   0,  -2,  -1,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   0,   1,   1,  -3,   4,   0,  -2,
   1,   3,   0,   0,   0,   0,  -1,   0,
   1,   0,   1,   1,   1,   0,   0,   0,
   0,   0,   0,   0,  -1,   0,   0,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  52,   0,   0,  -3,   5,   6,  -3,   3,
   3,  -4,   0,   2,   2,  -2,  -1,   0,
   1,  -1,   1,   0,  -1,   1,   0,  -1,
  -1,   1,   0,   0,   0,   0,   0,   0,
  -1,   1,   0,   0,   0,   0,  -1,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -3,   0,   2,   2,   3,   1,   1,
   0,   0,   1,   0,  -1,   0,   1,   0,
   0,   0,  -1,   0,   1,   0,   0,   0,
   0,   0,   0,   1,   0,   0,   0,   1,
   0,   0,   1,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  40, -26,   6,   7,   6, -22,  -6,   0,
   2,  -3,   0,  -4,   2,  -3,  -2,  -2,
  -3,  -1,  -2,   0,   3,  -1,   3,   0,
   2,  -1,   0,  -1,  -1,   0,  -1,   1,
   0,   0,  -1,   0,  -1,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   3,   0,   1,  -3,   1,  -1,   2,
  -1,  -1,   0,  -1,  -1,  -2,  -1,   1,
   0,   1,   0,   1,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,  -4,   0,   0,   2,   2,  -2,   1,
  -1,  -4,   2,  -1,   1,   0,  -1,   0,
   0,   0,   1,   0,   1,   1,   1,  -1,
   0,   0,   0,   1,   0,   0,   0,   0,
   0,   0,   0,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,   0,   2,   5,   3,  -2,   3,   1,
   2,  -1,  -2,  -3,  -2,  -2,   1,   0,
   0,  -1,   2,  -1,   2,   0,   1,   1,
   1,   0,  -1,   0,   0,   0,   1,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,  -2,   3,   0,   1,  -1,  -2,   0,
   0,   3,  -1,   1,   0,   3,   0,   0,
   1,  -1,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,   0,  -1,  -1,  -2,   1,   1,   0,
   0,   1,  -1,   0,   0,   0,   0,   0,
   0,   1,   0,   1,   0,   0,  -1,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,  -1,  -3,   0,  -1,   3,   0,   1,
   0,   0,   1,  -1,  -1,   0,  -1,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   1,  -1,  -1,  -2,   4,  -1,   1,
  -1,  -2,   0,   1,   1,   1,   1,  -1,
   0,   1,   1,  -1,   0,  -1,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   0,  -1,   0,   1,   2,   2,   0,
   0,  -3,   1,   0,   1,  -1,   1,   0,
   0,  -1,   1,   1,   1,   0,   0,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,  -1,  -1,   2,   1,   1,  -1,   1,
   1,   1,   1,   0,  -1,   0,   0,   0,
   0,   0,  -1,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   1,   0,   0,   1,  -2,   0,   2,
   1,   0,   1,   0,  -1,   0,   0,   0,
   0,  -1,   0,   0,   0,   0,   1,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,  -1,   1,  -1,  -1,  -2,   1,  -1,
   0,  -1,   1,   1,  -1,  -1,  -1,   0,
   0,   0,   0,   0,  -1,  -1,   0,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,   0,   0,   0,  -4,  -7,  -3,   1,
   4,   2,  -2,   0,   0,   0,   1,  -1,
   0,   0,   2,  -1,  -1,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,  -1,   4,   1,   0,   6,   0,  -2,
  -1,   1,   1,   0,   0,   0,  -1,   0,
   0,   0,  -1,   1,  -4,   1,   0,   0,
   1,   1,   0,   0,   0,   0,   0,   1,
   0,   1,   0,   0,   0,  -1,   0,  -1,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,  -3,   1,  -4,   0,   2,   0,   1,
  -2,   0,  -1,   1,   3,   0,  -1,   0,
  -1,   0,   0,  -1,   0,   0,   0,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -2,   3,   3,   1,   2,   3,  -1,
   1,  -1,   1,  -1,  -1,   0,   1,   0,
   1,   0,   0,   2,   0,   0,  -1,   0,
   0,   0,   0,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  40, -16,  -4,  -3,   4, -24, -13,  -1,
  -2,   1,   1,  -3,  -2,  -1,  -6,  -2,
   0,   0,   2,   1,   1,   1,  -1,   1,
  -1,   0,  -1,  -1,  -1,   0,   0,   0,
   0,   0,   0,   1,  -1,   1,   0,   0,
   0,   0,   0,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,   5,  -2,  -1,  -1,   0,   0,   0,
   0,  -1,  -2,   1,  -2,   0,  -1,   0,
   0,   0,   1,   1,   1,  -1,   0,   1,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,  -3,   2,  -1,  -3,  -1,  -3,  -1,
   1,   3,  -1,   0,  -1,   1,  -1,   0,
   0,   0,  -1,   0,   0,   0,   0,   1,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -3,   0,   2,   0,  -4,   6,  -1,
   1,   0,  -2,   2,   0,   0,   1,   1,
   0,  -1,   0,   1,  -1,   1,  -1,  -1,
   1,  -1,   0,  -1,   0,   0,   0,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,  -7,   0,   0,  -1,  -7,  -4,  -1,
  -1,   0,  -1,   1,   0,  -2,  -2,  -1,
   0,   0,   0,  -1,   0,   0,   1,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   3,   0,   2,   0,  -1,   1,   2,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,  -1,   0,  -2,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   0,  -1,  -1,   2,   1,   0,  -2,
   1,  -1,  -4,   1,   0,   0,   0,   0,
   0,   0,  -1,   0,  -1,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,   2,  -1,  -1,   1,   0,  -2,   0,
   0,  -2,  -1,   0,   0,  -1,   1,   0,
   1,  -1,   0,   0,   0,   0,  -1,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   2,  -1,   0,  -2,   0,   0,   1,
  -1,   0,   0,   0,   0,   0,   2,   0,
   1,   1,   0,  -1,  -1,   1,   1,   0,
   0,   0,   0,  -1,   0,  -1,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,   0,  -2,  -1,   1,  -1,  -1,   1,
  -1,  -1,  -1,  -1,   0,   0,   0,   0,
   0,   0,   0,   1,  -1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   0,   0,   0,   1,   0,   1,   0,
   2,   0,   0,   0,   1,   0,   0,   0,
   0,   0,   0,  -1,   0,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   4,  -2,  -1,   0,  -6,   2,  -2,
   1,   3,   1,   0,   0,   1,  -2,   1,
   0,   1,   2,   1,  -1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -7,   6,   3,   6, -10,  -3,   3,
  -2,   1,  -2,   1,   3,   1,  -1,  -1,
   1,   1,  -1,   1,   1,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,  -1,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,   1,   2,  -2,   5,   3,   1,  -4,
   0,   5,  -2,   1,   1,   0,   0,   1,
  -1,   1,  -2,  -1,   0,  -1,   1,   0,
  -1,   1,   0,   0,  -1,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  53,  -4,  -5,  -3,  -2,   5,   1,   0,
  -2,   0,  -3,  -1,   3,   1,  -1,   0,
  -1,   2,   0,   0,  -2,  -1,  -1,   1,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,  -2,  -2,   0,  -4,   3,   1,  -1,
   0,   1,   0,   0,   1,   1,   1,   0,
   1,   0,   0,   1,   0,   1,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  38, -18,   7,  -3,   1, -19, -13,   1,
   2,  -5,   3,   1,   2,  -1,  -3,  -3,
  -2,   2,   0,   1,  -3,   2,   0,   0,
   0,   0,   0,  -1,   0,   0,  -1,   0,
   0,   0,   1,  -1,   0,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,   3,   0,   3,   2,   3,   2,   0,
  -2,  -1,  -1,   0,   0,   1,  -1,   0,
   1,   0,   0,  -1,   1,   0,  -1,   1,
   0,   0,   0,   0,   0,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  52,  -5,  -7,  -1,  -3,   9,   0,   2,
   0,  -2,  -3,   0,   0,   0,  -3,   0,
  -1,  -1,   1,  -1,   1,   0,   2,   2,
   1,   0,   0,   1,   0,   1,   0,   0,
   0,   1,   1,   0,   0,   0,   0,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,   1,  -5,  -1,  -1,   5,   5,   3,
   0,   0,   0,  -1,  -2,   2,  -1,   0,
   0,   1,   0,  -1,   2,   0,  -1,   1,
   0,   0,   0,  -1,  -1,   0,   0,   1,
   0,   0,   0,   1,   0,  -1,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,  -5,   0,   1,   3,  -6,  -2,   3,
  -1,   3,   1,   1,   0,   2,  -1,  -1,
   1,  -1,   0,   1,   1,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,   1,   3,   0,   0,   4,   0,  -1,
   1,   0,   0,  -1,   1,   0,   0,  -1,
   1,   0,   0,   1,  -1,   0,   0,   0,
   0,   0,   0,   0,   1,   0,   0,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  62,   0,   0,   1,   0,   1,   0,   0,
   0,  -1,  -1,   1,   0,   0,   0,   0,
   0,   0,   1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   0,   2,   4,   1,   0,   0,   1,
   2,  -1,   0,  -3,  -1,   0,   2,   0,
   0,   0,   0,   1,   1,  -1,   0,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   2,  -1,   0,  -1,   1,   0,   2,
  -2,  -1,   0,   1,   1,   1,   1,   0,
   0,   0,   0,   0,  -1,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,   0,   0,   2,   1,   0,  -1,  -1,
   0,  -1,   0,   0,  -1,   0,   0,   0,
   0,   1,   0,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   1,  -2,   3,   0,   2,  -1,   0,
   0,   0,  -2,   0,  -2,  -1,  -1,   0,
   0,   1,   0,   0,  -2,   0,   0,   1,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,  -1,  -2,   0,   1,  -2,   1,   0,
  -1,  -1,   2,  -1,   0,   0,   0,   0,
   0,  -1,  -1,   1,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,  -2,  -3,   1,  -1,  -4,  -4,   0,
  -7,   1,   0,  -1,  -2,  -1,   1,   0,
   1,   1,  -1,   2,   0,   0,   1,   0,
   0,  -1,   0,   0,   0,   0,   1,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   3,   0,   2,   1,   3,  -1,  -1,
  -1,  -2,   0,   0,  -1,   1,   0,   1,
   0,   1,   0,  -1,   1,   0,   0,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -2,   1,   2,   1,  -3,  -2,   0,
   3,  -4,   1,  -1,  -1,   0,  -1,   0,
   0,   1,  -2,   1,   0,   0,   1,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   1,   1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  50,  -1,   3,   1,   1,  11,   2,   2,
   0,  -3,   2,  -1,  -1,  -2,  -1,   0,
  -2,  -1,   0,   0,  -1,   1,   0,  -1,
   0,   0,   0,   1,  -1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  38, -20,  -1,  -1,  -3, -27, -14,   1,
  -1,  -1,   2,   4,   0,  -2,  -4,  -3,
   0,  -1,   1,   4,   0,   0,   0,   2,
   1,   1,   0,   1,  -1,  -1,   0,   0,
   0,   1,   0,  -1,   0,   0,   0,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,   3,   3,   0,   0,   3,   0,  -2,
   0,  -1,   1,   1,   2,   0,  -1,   0,
   1,   0,  -1,   1,   1,   0,  -1,   1,
   1,   0,   0,   0,  -1,   0,   0,   0,
  -1,   0,   0,   0,   0,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -6,  -1,  -1,   1,  -2,  -1,  -1,
  -2,  -1,   0,   0,  -1,  -2,   0,   0,
   0,  -2,   1,   0,   0,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,  -1,   2,   4,  -1,  -1,   4,   0,
   2,   1,  -1,   1,   0,  -2,   1,   0,
   0,   0,   0,   0,  -1,   0,   0,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,  -3,   0,  -1,   1,  -3,  -2,   1,
  -1,   2,   2,   0,  -1,  -1,  -1,   0,
   0,   0,   1,   1,   0,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,   2,   1,   0,   0,   5,   1,   0,
   1,   1,   0,   0,  -2,   1,  -1,   0,
   0,   1,   0,   0,   1,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   1,   0,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,  -1,   0,  -2,   2,   0,   0,  -1,
  -2,   0,  -1,  -1,   0,   0,   1,   0,
   0,   0,   0,   0,  -1,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,  -2,  -2,   3,   0,   1,   1,   0,
   4,   0,  -1,   1,   1,   1,   1,   0,
   0,   0,   0,  -2,  -1,   0,  -1,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   3,   0,   0,   0,  -1,   1,  -1,
  -4,  -1,   1,   1,   1,   0,   0,   0,
  -1,   0,   0,   0,   0,   0,   1,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,  -1,  -1,   1,  -1,   1,  -1,   0,
   1,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   2,   0,   1,   0,  -1,   1,   1,
   1,   1,   0,   0,   0,   0,   0,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,  -1,   1,   2,   2,  -5,   1,   0,
  -2,   0,   1,  -1,   1,  -1,  -1,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,  -6,   4,   1,   5,  -6,  -2,   2,
   2,  -2,   1,  -2,   2,   0,   1,   0,
   0,   0,  -1,   1,   0,   0,  -1,   1,
   0,   0,   0,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,   2,   0,  -1,  -3,   2,   2,   3,
   0,  -1,   2,   0,   1,   0,  -1,   0,
  -1,   0,   0,   0,  -1,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   1,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,  -2,   4,   0,   2,   2,  -4,   0,
   1,   1,   2,   0,   2,   1,  -1,   0,
   1,   1,  -1,   0,   1,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   1,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   1,  -3,  -3,  -2,   1,   1,   0,
  -1,  -4,   0,   0,   1,   2,   1,  -1,
   0,   1,   1,  -1,   1,   0,  -1,   1,
   1,   0,   0,   1,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  40, -25,   3,  -3,  -5, -19, -12,  -1,
  -1,   1,   2,   2,  -4,   4,  -4,  -1,
   2,   0,   1,   0,   2,   1,   2,  -1,
   1,   1,   0,  -1,  -1,   0,   0,   0,
   0,   1,   0,   0,   1,   0,  -1,  -1,
   0,   0,   0,   0,   0,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  52,   5,   5,   2,  -1,   5,  -3,  -3,
  -1,  -4,   3,   0,  -1,   1,   1,  -1,
   0,   0,   4,   1,  -1,   0,   2,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   1,   0,   0,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,  -3,   2,   0,   2,  -2,  -2,   0,
   1,   1,   3,  -2,   0,   0,  -1,   0,
   0,   0,   0,   1,   0,   0,   0,   1,
  -1,   0,   0,   0,  -1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  56,   1,  -3,   0,  -1,  -3,   4,   1,
   2,   1,  -1,  -1,  -3,   1,   0,   1,
   1,   0,   1,   1,   2,   0,   0,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   1,   0,   0,   0,   0,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,  -6,  -2,   1,  -1,  -6,  -3,  -2,
   0,  -1,  -1,  -2,   0,  -1,  -1,  -1,
  -1,   0,  -1,  -2,   0,   0,   0,  -1,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   3,   0,   0,  -2,   0,   0,  -1,
   1,   0,   1,   0,  -1,   0,   0,   0,
   0,   0,   2,   0,   2,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,   0,   2,   1,   0,   2,   0,   0,
   0,  -3,   0,   0,   0,   0,   0,   0,
   0,   0,   1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   2,   1,   0,   1,   1,   0,  -1,
  -1,   2,  -1,   0,   0,   0,   1,  -1,
   0,   1,  -1,   0,   1,   0,   0,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   2,   1,   1,  -1,   0,   1,  -1,
  -1,   1,   0,  -2,   0,   0,   0,   0,
  -1,   0,   2,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,  -1,   1,   1,   1,   2,  -2,   1,
   1,   0,   0,   1,  -1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,  -3,  -1,  -2,   0,  -1,  -1,  -1,
  -2,   0,   1,   1,   1,  -1,  -1,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,  -3,   0,   0,   1,  -2,   0,  -1,
   1,   1,  -2,   2,   0,   1,  -1,   0,
   0,   0,  -1,  -1,   0,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  51,  -7,   5,   0,   2, -14,  -4,   5,
   2,   1,  -1,   0,  -1,   0,   1,   0,
   0,   0,   0,  -1,   0,   0,   1,   0,
   0,   0,   0,   1,   0,   0,   0,   0,
   0,   0,  -1,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   0,   2,  -1,   0,   2,   0,   0,
   0,   0,   1,   1,  -2,   0,  -1,   1,
   0,   0,  -1,   0,   0,   0,   1,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  46,  -4,   6,  -4,   0,   5,  -2,  -4,
  -4,  -8,   3,   4,   0,   2,   2,   1,
   0,   0,   2,  -2,  -3,   0,  -1,  -2,
  -1,   0,   0,   0,   0,   0,   1,   1,
   0,   1,   1,   0,   0,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  53,  -6,   0,   1,  -1,   9,   4,  -3,
   0,   0,   0,  -1,   0,   0,   0,   0,
   1,   0,   1,   0,   1,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,  -1,   0,  -1,  -1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  36, -23,  -1,  -5,   5, -24, -11,   0,
  -4,   4,   2,   0,  -1,   2,  -3,  -2,
   0,   1,   1,   4,   2,   0,   3,  -3,
   1,   1,   1,   0,  -1,   0,   0,  -1,
   0,   0,   1,   1,   0,   0,   0,   0,
   0,   0,  -1,   0,  -1,   0,  -1,  -1,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,   6,  -2,   2,   0,  -2,   2,  -2,
  -3,   0,  -2,  -1,   1,   1,  -3,   1,
   1,   0,   1,   0,   1,   0,  -1,   0,
   0,   0,  -1,   0,   0,   0,  -1,   0,
   0,   1,   0,   0,   0,   0,   0,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  52,  -8,   0,   3,   0,  -2,  -4,  -1,
   3,  -2,   0,  -1,   3,   1,  -3,   0,
   2,   1,   1,  -2,  -2,   0,   0,  -1,
  -1,   1,   0,   1,   0,   0,   0,  -1,
   0,   0,   1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   1,   0,   1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -1,  -2,  -1,   1,  -2,   6,  -3,
   0,   1,   1,  -1,  -2,   0,   0,   0,
  -1,   1,   0,   0,   0,   0,   0,   1,
   0,   1,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   0,  -3,   1,   0,  -2,  -3,  -2,
   1,   2,   0,   2,   2,  -2,  -1,   0,
  -1,   0,   1,   1,  -2,   0,   0,   0,
   1,   0,   0,  -1,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   1,   1,   0,   1,   1,   1,  -3,
   1,   0,   1,   1,   1,  -1,   0,   0,
   0,   0,   0,   0,  -1,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
  -1,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,  -1,  -2,  -1,   0,   0,   0,   1,
   1,  -1,   0,   0,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   2,  -1,   3,  -1,   1,   0,   1,
  -4,   0,  -1,   1,   0,   1,   2,  -1,
   0,   1,  -1,   1,   0,   0,  -1,   0,
  -1,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,   0,   0,   0,   1,   1,   0,  -1,
   1,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,  -1,   0,   0,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,   1,   0,   1,   0,   2,   0,  -1,
   0,   1,   0,   0,   0,   1,   0,   0,
   1,   0,   0,   0,  -2,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,   0,  -2,   0,  -1,   1,   0,   1,
   0,  -2,   0,  -1,   2,   1,   1,   0,
   0,   0,   1,  -1,   0,   0,   0,   0,
   1,   0,   0,  -1,   0,   0,   0,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   1,  -2,   1,  -1,  -1,   2,   2,
   2,  -1,  -1,   0,  -2,   1,  -3,   0,
   0,   1,  -2,   1,   0,   0,   0,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   1,   0,   0,   0,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -7,   1,  -1,   0, -11,  -4,   1,
  -4,  -1,  -3,  -3,  -2,   2,  -1,  -1,
   1,  -1,  -1,  -3,  -2,  -1,  -1,  -1,
  -1,   0,   1,   0,   0,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   0,   3,   0,   4,   3,   0,  -2,
   0,   0,   0,  -2,   1,  -1,  -1,   0,
   0,   0,   1,   1,  -2,   0,   0,  -1,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  53,  -7,  -4,   3,  -3,   1,   0,   0,
   5,  -1,  -2,   1,   0,   0,   1,   0,
   0,   0,   1,   0,  -2,   0,   0,   1,
   1,   1,   0,   0,   0,   0,   0,   1,
   0,   0,   0,   0,   1,   0,   0,   0,
   0,  -1,   0,   0,  -1,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  52,   2,   1,  -1,  -4,   3,   2,   3,
   3,   2,   2,  -1,  -2,  -1,   0,   0,
   0,   0,  -1,  -1,   1,  -1,  -2,  -1,
  -1,   0,   1,   0,  -1,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  40, -24,  -4,   0,  -9, -20, -13,  -2,
   0,   0,   4,   3,  -1,   2,  -4,  -2,
   1,   2,   1,   0,   2,   1,   2,   0,
   0,   1,   1,   0,  -1,   0,   0,   0,
   0,   0,   2,   1,   1,   1,  -1,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,   2,   0,  -3,  -3,   4,   0,   0,
  -2,  -2,   2,   0,   2,   1,  -2,   0,
   0,   0,   0,   0,  -1,   1,   1,  -1,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  53,  -6,   1,  -1,  -1,  -1,  -3,   2,
  -4,  -1,  -1,   0,  -2,   2,  -1,  -1,
  -1,  -1,  -1,  -1,  -2,  -1,  -1,   0,
  -2,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,  -1,   0,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,

  57,  -6,   0,  -4,   0,   0,   6,   2,
  -2,   0,  -1,   1,  -2,   0,   3,   1,
   0,   2,   0,   0,  -1,   0,  -1,   0,
   0,   1,   0,   0,   0,   0,   1,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,  -3,   1,  -2,   2,  -3,  -3,   2,
  -1,  -3,   1,  -2,  -2,   2,  -1,   0,
   1,   0,  -1,   0,   0,   0,  -1,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
   1,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   2,  -1,   1,  -1,  -1,   1,   1,
  -1,  -1,   1,   0,   2,  -1,   0,   0,
   0,   0,   1,   0,  -1,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,  -2,  -2,   1,  -1,   1,   0,   0,
  -1,   2,   0,   0,  -1,   1,   0,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,   1,   0,  -1,  -1,   2,  -1,  -1,
   2,   1,   0,   0,   0,   0,   1,   0,
   0,  -2,  -1,   0,   0,   0,  -1,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,   2,   0,  -2,   0,   0,   1,  -1,
   0,   0,   0,   0,   1,   0,   1,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,   0,  -1,  -1,  -1,   1,  -2,  -1,
  -1,   1,   0,   0,   0,  -1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,  -1,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   3,   1,  -1,  -2,   3,  -1,  -1,
   0,  -3,   1,   1,   0,   1,   0,   0,
   0,  -1,   1,  -1,  -1,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,  -2,  -1,   0,   0,  -3,   2,   0,
   0,  -1,  -1,   0,  -1,   1,  -1,   0,
   0,  -1,   0,  -1,   0,   0,   0,   0,
   1,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  53,   0,   1,  -3,   5, -11,  -4,   4,
  -2,  -1,  -1,   0,  -2,   0,   1,  -1,
   2,  -2,   0,  -2,   0,   0,   0,   0,
  -1,   0,   0,   0,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,   6,  -2,  -1,  -1,   1,  -1,   3,
   2,   2,  -1,   1,   0,   0,   0,   0,
   0,   0,   0,   0,  -1,  -2,   0,   0,
   1,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  50,  -5,   2,  -3,   5,   4,  -3,   2,
   0,  -1,   3,  -3,  -2,  -2,   0,   1,
   1,  -2,  -2,   0,   1,   1,  -2,   0,
   1,   0,   0,   0,  -1,   0,   0,   1,
   1,   0,   0,   0,   0,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  51,   0,  -4,  -1,   4,  12,   1,   2,
   3,  -5,   1,  -1,   0,  -2,  -2,   0,
   0,  -2,   2,   3,   2,   0,   2,  -1,
   0,   0,   0,   1,  -1,   0,   0,   1,
  -1,  -1,   0,   0,   0,   0,  -1,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  28, -28,   3,   5,  -7, -25, -11,   3,
   4,   3,  -4,   3,  -5,   2,  -2,  -2,
   1,  -3,   1,  -1,   2,  -2,  -2,  -1,
  -2,  -3,   0,   0,  -1,   0,  -2,  -1,
   1,   0,   0,   0,   0,   0,   0,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  52,   5,   0,   2,   1,   1,  -1,   3,
  -2,  -2,  -1,   2,  -3,   1,  -1,   0,
   0,   0,   0,   0,   0,   1,   2,   0,
   0,   0,   0,   0,  -1,   0,   0,   1,
  -1,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   1,

  53,  -5,   0,   0,   0,  -3,  -2,   1,
  -2,   1,   1,   4,  -4,   1,  -1,  -1,
   0,  -1,   1,  -1,   0,  -1,   0,  -2,
   0,   0,   0,   0,   0,   1,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,  -2,   0,   2,   1,  -3,   4,   0,
  -1,   0,  -3,  -2,   3,   0,   1,   0,
   0,   0,   0,  -1,   0,   0,   1,   0,
  -1,   0,   0,   0,  -1,   0,   0,   1,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,  -5,  -2,   0,  -1,  -5,  -1,  -1,
   1,   1,   1,   2,  -1,   0,  -1,   0,
   0,   0,   0,   1,   0,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   2,  -1,   2,   1,   0,   1,   0,
   0,  -2,   0,   0,  -1,   0,   1,   0,
   0,  -1,   0,   1,   2,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,  -1,  -1,  -1,  -1,   0,  -1,   0,
   1,   0,  -1,  -1,   0,  -1,   0,   0,
   0,   0,  -1,   0,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,  -1,  -1,  -1,   0,   2,   1,   1,
  -1,   1,   2,   1,   0,   1,   0,   0,
   0,   0,   0,   0,   1,   0,   0,  -1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,   3,  -1,  -1,   1,   0,   0,   0,
   1,  -1,   2,   1,  -1,  -1,   1,   0,
   0,   0,   0,  -1,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  60,  -2,   1,   0,   0,   1,   0,   1,
  -1,  -1,   1,   0,  -1,   1,   0,   0,
   0,   0,   0,   1,   1,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   3,  -2,   0,   1,   1,  -2,   1,
   1,  -1,  -2,   0,   2,   0,   0,   0,
   0,   0,   0,   0,  -1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,  -1,  -2,  -1,  -1,  -5,   2,  -1,
  -3,   1,  -1,  -2,   0,   0,  -1,   1,
   0,   0,   0,   0,   0,   0,  -1,  -1,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,  -1,   0,   2,   1,  -8,  -1,   1,
  -2,  -3,  -1,   0,   2,  -1,   0,   0,
   0,  -1,  -1,   1,   1,   0,  -1,   1,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,  -1,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,   1,   1,   2,  -2,   0,   2,   0,
   1,   0,  -1,  -1,   0,  -1,  -1,   0,
   0,   0,   0,   0,   1,   0,   1,   1,
   0,   0,   0,   0,  -1,   0,   0,   0,
   0,  -1,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,  -4,   0,   1,   0,   2,  -2,   1,
   0,   1,   0,   2,   0,   0,   0,   1,
  -1,   0,   1,   0,   1,   0,  -2,   1,
   1,   0,   0,   0,   0,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  51,  -2,   6,   3,   3,   6,   3,  -2,
   0,  -2,   0,  -1,   0,  -3,   0,   1,
  -1,  -1,   1,  -1,   0,   0,   1,   0,
  -1,   0,  -1,   1,  -1,  -1,   0,   0,
   0,   0,   0,   1,   0,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  37, -25,   8,  -6,   6, -22, -10,   3,
  -4,   6,   4,   1,  -2,  -5,  -3,  -1,
  -4,   3,   1,   2,  -1,   1,  -3,   0,
  -1,   1,  -1,   0,  -1,   0,   1,   0,
   1,   0,   1,  -1,  -1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  52,   5,   4,  -2,  -1,   2,  -1,  -3,
  -2,  -5,   1,   2,   1,   0,  -1,   0,
  -1,   0,  -1,  -2,   3,  -1,  -1,   1,
   0,   0,   1,   0,   0,   0,   0,   0,
   0,   0,   1,   1,   0,   0,   0,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  53,  -7,   3,  -1,   1,   0,  -2,  -1,
   0,   4,   1,   0,   0,   1,  -1,   0,
   0,   0,  -2,   1,   1,  -1,   0,   0,
   0,   1,   0,   1,   0,   0,   0,   0,
   0,   0,   1,   0,   0,   1,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,  -2,  -2,   1,   0,  -1,   5,  -2,
   2,   0,   0,   1,  -1,   0,   1,   1,
   1,  -1,   0,   0,  -1,   0,  -2,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  57,  -6,  -3,  -3,  -4,  -8,  -3,  -2,
  -1,  -1,  -1,  -2,   0,  -1,  -2,   0,
  -1,   0,  -1,   0,   1,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,  -1,   1,   1,  -1,   0,   0,   0,
   2,   1,  -2,   1,   0,   1,   0,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  62,   0,  -1,   0,   0,   1,   0,   1,
   0,   0,  -1,   0,   1,   0,   0,   0,
   0,   0,   1,   0,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  62,   1,   0,  -1,   0,   1,   0,   0,
   1,   0,   1,   0,   0,   0,   1,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  62,   0,  -1,  -1,   0,   0,   1,   0,
  -1,  -1,   0,   0,   1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,  -1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  61,   0,   0,   0,   1,   1,  -1,   0,
  -1,   3,  -1,   0,   2,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   1,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  59,   1,   1,  -2,   0,   1,   0,  -1,
   0,   0,  -2,  -1,  -1,   0,   0,   0,
   0,   0,   1,   0,  -1,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  55,   6,   0,  -4,   0, -11,   2,   0,
   2,   3,  -2,  -1,  -1,   0,  -3,   1,
  -1,   0,   2,   1,   1,   0,  -1,  -1,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,  -1,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,  -6,   2,  -3,   1,  -7,  -3,  -3,
   0,  -4,  -2,  -2,  -2,   0,   0,   0,
   0,   0,  -2,  -2,   1,   0,   1,   0,
  -1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,  -1,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  58,   0,   0,   0,   0,   2,   1,  -1,
  -2,   0,   0,   0,   0,   0,   0,   1,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,  -1,   2,  -1,  -3,   4,  -4,  -1,
   1,   3,  -1,  -1,   1,   2,  -1,   1,
   0,  -1,  -2,   1,   2,   0,   0,   1,
   0,   0,   0,   0,  -1,   1,   0,   0,
   0,  -1,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,

  54,   1,   5,  -2,   0,   5,   1,   0,
   0,   2,  -2,   0,  -1,  -1,  -1,   0,
  -1,   2,   1,  -1,   1,   0,  -1,   1,
  -1,   1,   0,   0,  -1,   0,   0,   0,
   1,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,   0,
   0,   0,   0,   0,   0,   0,   0,  -1  };

endmodule
