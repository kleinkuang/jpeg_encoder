// File:    ac_lut.py
// Author:  Lei Kuang
// Date:    13th July 2020
// @ Imperial College London

// Note that the actual length is len + 1
// e.g., len=4'd3 -> bin[3:0] are valid;

module ac_lut
(
    input  logic [3:0]  rrrr,
    input  logic [3:0]  ssss,
    output logic [4:0]  len,
    output logic [15:0] bin
);

logic [7:0] rrrrssss;

assign rrrrssss = {rrrr, ssss};

always_comb begin
    len = '0;
    case(rrrrssss)
        8'h00:   len = 5'd4;
        8'h01:   len = 5'd2;
        8'h02:   len = 5'd2;
        8'h03:   len = 5'd3;
        8'h04:   len = 5'd4;
        8'h05:   len = 5'd5;
        8'h06:   len = 5'd7;
        8'h07:   len = 5'd8;
        8'h08:   len = 5'd10;
        8'h09:   len = 5'd16;
        8'h0A:   len = 5'd16;

        8'h11:   len = 5'd4;
        8'h12:   len = 5'd5;
        8'h13:   len = 5'd7;
        8'h14:   len = 5'd9;
        8'h15:   len = 5'd11;
        8'h16:   len = 5'd16;
        8'h17:   len = 5'd16;
        8'h18:   len = 5'd16;
        8'h19:   len = 5'd16;
        8'h1A:   len = 5'd16;

        8'h21:   len = 5'd5;
        8'h22:   len = 5'd8;
        8'h23:   len = 5'd10;
        8'h24:   len = 5'd12;
        8'h25:   len = 5'd16;
        8'h26:   len = 5'd16;
        8'h27:   len = 5'd16;
        8'h28:   len = 5'd16;
        8'h29:   len = 5'd16;
        8'h2A:   len = 5'd16;

        8'h31:   len = 5'd6;
        8'h32:   len = 5'd9;
        8'h33:   len = 5'd12;
        8'h34:   len = 5'd16;
        8'h35:   len = 5'd16;
        8'h36:   len = 5'd16;
        8'h37:   len = 5'd16;
        8'h38:   len = 5'd16;
        8'h39:   len = 5'd16;
        8'h3A:   len = 5'd16;

        8'h41:   len = 5'd6;
        8'h42:   len = 5'd10;
        8'h43:   len = 5'd16;
        8'h44:   len = 5'd16;
        8'h45:   len = 5'd16;
        8'h46:   len = 5'd16;
        8'h47:   len = 5'd16;
        8'h48:   len = 5'd16;
        8'h49:   len = 5'd16;
        8'h4A:   len = 5'd16;

        8'h51:   len = 5'd7;
        8'h52:   len = 5'd11;
        8'h53:   len = 5'd16;
        8'h54:   len = 5'd16;
        8'h55:   len = 5'd16;
        8'h56:   len = 5'd16;
        8'h57:   len = 5'd16;
        8'h58:   len = 5'd16;
        8'h59:   len = 5'd16;
        8'h5A:   len = 5'd16;

        8'h61:   len = 5'd7;
        8'h62:   len = 5'd12;
        8'h63:   len = 5'd16;
        8'h64:   len = 5'd16;
        8'h65:   len = 5'd16;
        8'h66:   len = 5'd16;
        8'h67:   len = 5'd16;
        8'h68:   len = 5'd16;
        8'h69:   len = 5'd16;
        8'h6A:   len = 5'd16;

        8'h71:   len = 5'd8;
        8'h72:   len = 5'd12;
        8'h73:   len = 5'd16;
        8'h74:   len = 5'd16;
        8'h75:   len = 5'd16;
        8'h76:   len = 5'd16;
        8'h77:   len = 5'd16;
        8'h78:   len = 5'd16;
        8'h79:   len = 5'd16;
        8'h7A:   len = 5'd16;

        8'h81:   len = 5'd9;
        8'h82:   len = 5'd15;
        8'h83:   len = 5'd16;
        8'h84:   len = 5'd16;
        8'h85:   len = 5'd16;
        8'h86:   len = 5'd16;
        8'h87:   len = 5'd16;
        8'h88:   len = 5'd16;
        8'h89:   len = 5'd16;
        8'h8A:   len = 5'd16;

        8'h91:   len = 5'd9;
        8'h92:   len = 5'd16;
        8'h93:   len = 5'd16;
        8'h94:   len = 5'd16;
        8'h95:   len = 5'd16;
        8'h96:   len = 5'd16;
        8'h97:   len = 5'd16;
        8'h98:   len = 5'd16;
        8'h99:   len = 5'd16;
        8'h9A:   len = 5'd16;

        8'hA1:   len = 5'd9;
        8'hA2:   len = 5'd16;
        8'hA3:   len = 5'd16;
        8'hA4:   len = 5'd16;
        8'hA5:   len = 5'd16;
        8'hA6:   len = 5'd16;
        8'hA7:   len = 5'd16;
        8'hA8:   len = 5'd16;
        8'hA9:   len = 5'd16;
        8'hAA:   len = 5'd16;

        8'hB1:   len = 5'd10;
        8'hB2:   len = 5'd16;
        8'hB3:   len = 5'd16;
        8'hB4:   len = 5'd16;
        8'hB5:   len = 5'd16;
        8'hB6:   len = 5'd16;
        8'hB7:   len = 5'd16;
        8'hB8:   len = 5'd16;
        8'hB9:   len = 5'd16;
        8'hBA:   len = 5'd16;

        8'hC1:   len = 5'd10;
        8'hC2:   len = 5'd16;
        8'hC3:   len = 5'd16;
        8'hC4:   len = 5'd16;
        8'hC5:   len = 5'd16;
        8'hC6:   len = 5'd16;
        8'hC7:   len = 5'd16;
        8'hC8:   len = 5'd16;
        8'hC9:   len = 5'd16;
        8'hCA:   len = 5'd16;

        8'hD1:   len = 5'd11;
        8'hD2:   len = 5'd16;
        8'hD3:   len = 5'd16;
        8'hD4:   len = 5'd16;
        8'hD5:   len = 5'd16;
        8'hD6:   len = 5'd16;
        8'hD7:   len = 5'd16;
        8'hD8:   len = 5'd16;
        8'hD9:   len = 5'd16;
        8'hDA:   len = 5'd16;

        8'hE1:   len = 5'd16;
        8'hE2:   len = 5'd16;
        8'hE3:   len = 5'd16;
        8'hE4:   len = 5'd16;
        8'hE5:   len = 5'd16;
        8'hE6:   len = 5'd16;
        8'hE7:   len = 5'd16;
        8'hE8:   len = 5'd16;
        8'hE9:   len = 5'd16;
        8'hEA:   len = 5'd16;

        8'hF0:   len = 5'd11;
        8'hF1:   len = 5'd16;
        8'hF2:   len = 5'd16;
        8'hF3:   len = 5'd16;
        8'hF4:   len = 5'd16;
        8'hF5:   len = 5'd16;
        8'hF6:   len = 5'd16;
        8'hF7:   len = 5'd16;
        8'hF8:   len = 5'd16;
        8'hF9:   len = 5'd16;
        8'hFA:   len = 5'd16;
    endcase
end

always_comb begin
    bin = '0;
    case(rrrrssss)
        8'h00:   bin = 16'b1010;
        8'h01:   bin = 16'b0;
        8'h02:   bin = 16'b1;
        8'h03:   bin = 16'b100;
        8'h04:   bin = 16'b1011;
        8'h05:   bin = 16'b11010;
        8'h06:   bin = 16'b1111000;
        8'h07:   bin = 16'b11111000;
        8'h08:   bin = 16'b1111110110;
        8'h09:   bin = 16'b1111111110000010;
        8'h0A:   bin = 16'b1111111110000011;
        
        8'h11:   bin = 16'b1100;
        8'h12:   bin = 16'b11011;
        8'h13:   bin = 16'b1111001;
        8'h14:   bin = 16'b111110110;
        8'h15:   bin = 16'b11111110110;
        8'h16:   bin = 16'b1111111110000100;
        8'h17:   bin = 16'b1111111110000101;
        8'h18:   bin = 16'b1111111110000110;
        8'h19:   bin = 16'b1111111110000111;
        8'h1A:   bin = 16'b1111111110001000;
        
        8'h21:   bin = 16'b11100;
        8'h22:   bin = 16'b11111001;
        8'h23:   bin = 16'b1111110111;
        8'h24:   bin = 16'b111111110100;
        8'h25:   bin = 16'b1111111110001001;
        8'h26:   bin = 16'b1111111110001010;
        8'h27:   bin = 16'b1111111110001011;
        8'h28:   bin = 16'b1111111110001100;
        8'h29:   bin = 16'b1111111110001101;
        8'h2A:   bin = 16'b1111111110001110;
        
        8'h31:   bin = 16'b111010;
        8'h32:   bin = 16'b111110111;
        8'h33:   bin = 16'b111111110101;
        8'h34:   bin = 16'b1111111110001111;
        8'h35:   bin = 16'b1111111110010000;
        8'h36:   bin = 16'b1111111110010001;
        8'h37:   bin = 16'b1111111110010010;
        8'h38:   bin = 16'b1111111110010011;
        8'h39:   bin = 16'b1111111110010100;
        8'h3A:   bin = 16'b1111111110010101;
        
        8'h41:   bin = 16'b111011;
        8'h42:   bin = 16'b1111111000;
        8'h43:   bin = 16'b1111111110010110;
        8'h44:   bin = 16'b1111111110010111;
        8'h45:   bin = 16'b1111111110011000;
        8'h46:   bin = 16'b1111111110011001;
        8'h47:   bin = 16'b1111111110011010;
        8'h48:   bin = 16'b1111111110011011;
        8'h49:   bin = 16'b1111111110011100;
        8'h4A:   bin = 16'b1111111110011101;
        
        8'h51:   bin = 16'b1111010;
        8'h52:   bin = 16'b11111110111;
        8'h53:   bin = 16'b1111111110011110;
        8'h54:   bin = 16'b1111111110011111;
        8'h55:   bin = 16'b1111111110100000;
        8'h56:   bin = 16'b1111111110100001;
        8'h57:   bin = 16'b1111111110100010;
        8'h58:   bin = 16'b1111111110100011;
        8'h59:   bin = 16'b1111111110100100;
        8'h5A:   bin = 16'b1111111110100101;
        
        8'h61:   bin = 16'b1111011;
        8'h62:   bin = 16'b111111110110;
        8'h63:   bin = 16'b1111111110100110;
        8'h64:   bin = 16'b1111111110100111;
        8'h65:   bin = 16'b1111111110101000;
        8'h66:   bin = 16'b1111111110101001;
        8'h67:   bin = 16'b1111111110101010;
        8'h68:   bin = 16'b1111111110101011;
        8'h69:   bin = 16'b1111111110101100;
        8'h6A:   bin = 16'b1111111110101101;
        
        8'h71:   bin = 16'b11111010;
        8'h72:   bin = 16'b111111110111;
        8'h73:   bin = 16'b1111111110101110;
        8'h74:   bin = 16'b1111111110101111;
        8'h75:   bin = 16'b1111111110110000;
        8'h76:   bin = 16'b1111111110110001;
        8'h77:   bin = 16'b1111111110110010;
        8'h78:   bin = 16'b1111111110110011;
        8'h79:   bin = 16'b1111111110110100;
        8'h7A:   bin = 16'b1111111110110101;
        
        8'h81:   bin = 16'b111111000;
        8'h82:   bin = 16'b111111111000000;
        8'h83:   bin = 16'b1111111110110110;
        8'h84:   bin = 16'b1111111110110111;
        8'h85:   bin = 16'b1111111110111000;
        8'h86:   bin = 16'b1111111110111001;
        8'h87:   bin = 16'b1111111110111010;
        8'h88:   bin = 16'b1111111110111011;
        8'h89:   bin = 16'b1111111110111100;
        8'h8A:   bin = 16'b1111111110111101;
        
        8'h91:   bin = 16'b111111001;
        8'h92:   bin = 16'b1111111110111110;
        8'h93:   bin = 16'b1111111110111111;
        8'h94:   bin = 16'b1111111111000000;
        8'h95:   bin = 16'b1111111111000001;
        8'h96:   bin = 16'b1111111111000010;
        8'h97:   bin = 16'b1111111111000011;
        8'h98:   bin = 16'b1111111111000100;
        8'h99:   bin = 16'b1111111111000101;
        8'h9A:   bin = 16'b1111111111000110;
        
        8'hA1:   bin = 16'b111111010;
        8'hA2:   bin = 16'b1111111111000111;
        8'hA3:   bin = 16'b1111111111001000;
        8'hA4:   bin = 16'b1111111111001001;
        8'hA5:   bin = 16'b1111111111001010;
        8'hA6:   bin = 16'b1111111111001011;
        8'hA7:   bin = 16'b1111111111001100;
        8'hA8:   bin = 16'b1111111111001101;
        8'hA9:   bin = 16'b1111111111001110;
        8'hAA:   bin = 16'b1111111111001111;
        
        8'hB1:   bin = 16'b1111111001;
        8'hB2:   bin = 16'b1111111111010000;
        8'hB3:   bin = 16'b1111111111010001;
        8'hB4:   bin = 16'b1111111111010010;
        8'hB5:   bin = 16'b1111111111010011;
        8'hB6:   bin = 16'b1111111111010100;
        8'hB7:   bin = 16'b1111111111010101;
        8'hB8:   bin = 16'b1111111111010110;
        8'hB9:   bin = 16'b1111111111010111;
        8'hBA:   bin = 16'b1111111111011000;
        
        8'hC1:   bin = 16'b1111111010;
        8'hC2:   bin = 16'b1111111111011001;
        8'hC3:   bin = 16'b1111111111011010;
        8'hC4:   bin = 16'b1111111111011011;
        8'hC5:   bin = 16'b1111111111011100;
        8'hC6:   bin = 16'b1111111111011101;
        8'hC7:   bin = 16'b1111111111011110;
        8'hC8:   bin = 16'b1111111111011111;
        8'hC9:   bin = 16'b1111111111100000;
        8'hCA:   bin = 16'b1111111111100001;
        
        8'hD1:   bin = 16'b11111111000;
        8'hD2:   bin = 16'b1111111111100010;
        8'hD3:   bin = 16'b1111111111100011;
        8'hD4:   bin = 16'b1111111111100100;
        8'hD5:   bin = 16'b1111111111100101;
        8'hD6:   bin = 16'b1111111111100110;
        8'hD7:   bin = 16'b1111111111100111;
        8'hD8:   bin = 16'b1111111111101000;
        8'hD9:   bin = 16'b1111111111101001;
        8'hDA:   bin = 16'b1111111111101010;
        
        8'hE1:   bin = 16'b1111111111101011;
        8'hE2:   bin = 16'b1111111111101100;
        8'hE3:   bin = 16'b1111111111101101;
        8'hE4:   bin = 16'b1111111111101110;
        8'hE5:   bin = 16'b1111111111101111;
        8'hE6:   bin = 16'b1111111111110000;
        8'hE7:   bin = 16'b1111111111110001;
        8'hE8:   bin = 16'b1111111111110010;
        8'hE9:   bin = 16'b1111111111110011;
        8'hEA:   bin = 16'b1111111111110100;
        
        8'hF0:   bin = 16'b11111111001;
        8'hF1:   bin = 16'b1111111111110101;
        8'hF2:   bin = 16'b1111111111110110;
        8'hF3:   bin = 16'b1111111111110111;
        8'hF4:   bin = 16'b1111111111111000;
        8'hF5:   bin = 16'b1111111111111001;
        8'hF6:   bin = 16'b1111111111111010;
        8'hF7:   bin = 16'b1111111111111011;
        8'hF8:   bin = 16'b1111111111111100;
        8'hF9:   bin = 16'b1111111111111101;
        8'hFA:   bin = 16'b1111111111111110;
        
    endcase
end

endmodule
