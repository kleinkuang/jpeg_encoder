// File:    fdct_tb.sv
// Author:  Lei Kuang
// Date:    17th June 2020
// @ Imperial College London

module fdct_tb;

logic        clk;
logic        nrst;
logic [7:0]  din;
logic        din_valid;
logic [7:0]  dout;
logic        dout_valid;

fdct dut(.*);

initial begin
    clk = '0;
    forever #5ns clk = ~clk;
end

logic [13:0] din_cnt;
logic [7:0]  img [16383:0];

initial begin
    nrst      = '0;
    din_cnt   = '0;
    din_valid = '0;
    
    @(posedge clk)
        nrst <= '1;
    
    forever begin
        @(posedge clk) begin
            din_valid <= ~din_valid;

            if(din_valid)
                din_cnt <= din_cnt + 1;
        end
    end
end

assign din = img[din_cnt];

initial begin
    byte temp;
    integer cnt = 0;
    
    forever @ (negedge clk) begin
        if(dout_valid) begin
            if(cnt % 64 == 0)
                 $write("MCU: %d\n", cnt >> 6);

            temp = dout;
            $write("%6d", temp);

            cnt = cnt + 1;
            if(cnt % 8 == 0)
                $write("\n");

        end
    end
end

// Debug
logic [5:0] pix_cnt;
logic [7:0] mcu_cnt;

logic end_of_mcu;
logic end_of_img;

assign end_of_mcu = pix_cnt=='1;
assign end_of_img = mcu_cnt=='1;

always_ff @ (posedge clk, negedge nrst)
    if(~nrst) begin
        pix_cnt <= '0;
        mcu_cnt <= '0;
    end
    else begin
        if(dout_valid)
            pix_cnt <= pix_cnt + 6'd1;
        if(end_of_mcu)
            mcu_cnt <= mcu_cnt + 8'd1; 
    end

// ROM Assignment
assign img[    0] = 255;
assign img[    1] = 255;
assign img[    2] = 255;
assign img[    3] = 255;
assign img[    4] = 255;
assign img[    5] = 255;
assign img[    6] = 255;
assign img[    7] = 255;
assign img[    8] = 255;
assign img[    9] = 255;
assign img[   10] = 255;
assign img[   11] = 255;
assign img[   12] = 255;
assign img[   13] = 255;
assign img[   14] = 255;
assign img[   15] = 255;
assign img[   16] = 255;
assign img[   17] = 255;
assign img[   18] = 255;
assign img[   19] = 255;
assign img[   20] = 255;
assign img[   21] = 255;
assign img[   22] = 255;
assign img[   23] = 255;
assign img[   24] = 255;
assign img[   25] = 255;
assign img[   26] = 255;
assign img[   27] = 255;
assign img[   28] = 255;
assign img[   29] = 255;
assign img[   30] = 255;
assign img[   31] = 255;
assign img[   32] = 255;
assign img[   33] = 255;
assign img[   34] = 255;
assign img[   35] = 255;
assign img[   36] = 255;
assign img[   37] = 255;
assign img[   38] = 255;
assign img[   39] = 255;
assign img[   40] = 255;
assign img[   41] = 255;
assign img[   42] = 255;
assign img[   43] = 255;
assign img[   44] = 255;
assign img[   45] = 255;
assign img[   46] = 255;
assign img[   47] = 255;
assign img[   48] = 255;
assign img[   49] = 255;
assign img[   50] = 255;
assign img[   51] = 255;
assign img[   52] = 255;
assign img[   53] = 255;
assign img[   54] = 255;
assign img[   55] = 255;
assign img[   56] = 255;
assign img[   57] = 255;
assign img[   58] = 255;
assign img[   59] = 255;
assign img[   60] = 255;
assign img[   61] = 255;
assign img[   62] = 255;
assign img[   63] = 255;
assign img[   64] = 255;
assign img[   65] = 255;
assign img[   66] = 255;
assign img[   67] = 255;
assign img[   68] = 255;
assign img[   69] = 255;
assign img[   70] = 255;
assign img[   71] = 255;
assign img[   72] = 255;
assign img[   73] = 255;
assign img[   74] = 255;
assign img[   75] = 255;
assign img[   76] = 255;
assign img[   77] = 255;
assign img[   78] = 255;
assign img[   79] = 255;
assign img[   80] = 255;
assign img[   81] = 255;
assign img[   82] = 255;
assign img[   83] = 255;
assign img[   84] = 255;
assign img[   85] = 255;
assign img[   86] = 255;
assign img[   87] = 255;
assign img[   88] = 255;
assign img[   89] = 255;
assign img[   90] = 255;
assign img[   91] = 255;
assign img[   92] = 255;
assign img[   93] = 255;
assign img[   94] = 255;
assign img[   95] = 255;
assign img[   96] = 255;
assign img[   97] = 255;
assign img[   98] = 255;
assign img[   99] = 255;
assign img[  100] = 255;
assign img[  101] = 255;
assign img[  102] = 255;
assign img[  103] = 255;
assign img[  104] = 255;
assign img[  105] = 255;
assign img[  106] = 255;
assign img[  107] = 255;
assign img[  108] = 255;
assign img[  109] = 255;
assign img[  110] = 255;
assign img[  111] = 255;
assign img[  112] = 255;
assign img[  113] = 255;
assign img[  114] = 255;
assign img[  115] = 255;
assign img[  116] = 255;
assign img[  117] = 255;
assign img[  118] = 255;
assign img[  119] = 255;
assign img[  120] = 255;
assign img[  121] = 255;
assign img[  122] = 255;
assign img[  123] = 255;
assign img[  124] = 255;
assign img[  125] = 255;
assign img[  126] = 255;
assign img[  127] = 255;
assign img[  128] = 255;
assign img[  129] = 255;
assign img[  130] = 255;
assign img[  131] = 255;
assign img[  132] = 255;
assign img[  133] = 255;
assign img[  134] = 255;
assign img[  135] = 255;
assign img[  136] = 255;
assign img[  137] = 255;
assign img[  138] = 255;
assign img[  139] = 255;
assign img[  140] = 255;
assign img[  141] = 255;
assign img[  142] = 255;
assign img[  143] = 255;
assign img[  144] = 255;
assign img[  145] = 255;
assign img[  146] = 255;
assign img[  147] = 255;
assign img[  148] = 255;
assign img[  149] = 255;
assign img[  150] = 255;
assign img[  151] = 255;
assign img[  152] = 255;
assign img[  153] = 255;
assign img[  154] = 255;
assign img[  155] = 255;
assign img[  156] = 255;
assign img[  157] = 255;
assign img[  158] = 255;
assign img[  159] = 255;
assign img[  160] = 255;
assign img[  161] = 255;
assign img[  162] = 255;
assign img[  163] = 255;
assign img[  164] = 255;
assign img[  165] = 255;
assign img[  166] = 255;
assign img[  167] = 255;
assign img[  168] = 255;
assign img[  169] = 255;
assign img[  170] = 255;
assign img[  171] = 255;
assign img[  172] = 255;
assign img[  173] = 255;
assign img[  174] = 255;
assign img[  175] = 255;
assign img[  176] = 255;
assign img[  177] = 255;
assign img[  178] = 255;
assign img[  179] = 255;
assign img[  180] = 255;
assign img[  181] = 255;
assign img[  182] = 255;
assign img[  183] = 255;
assign img[  184] = 255;
assign img[  185] = 255;
assign img[  186] = 255;
assign img[  187] = 255;
assign img[  188] = 255;
assign img[  189] = 255;
assign img[  190] = 255;
assign img[  191] = 255;
assign img[  192] = 255;
assign img[  193] = 255;
assign img[  194] = 255;
assign img[  195] = 255;
assign img[  196] = 255;
assign img[  197] = 255;
assign img[  198] = 255;
assign img[  199] = 255;
assign img[  200] = 255;
assign img[  201] = 255;
assign img[  202] = 255;
assign img[  203] = 255;
assign img[  204] = 255;
assign img[  205] = 255;
assign img[  206] = 255;
assign img[  207] = 255;
assign img[  208] = 255;
assign img[  209] = 255;
assign img[  210] = 255;
assign img[  211] = 255;
assign img[  212] = 255;
assign img[  213] = 255;
assign img[  214] = 255;
assign img[  215] = 255;
assign img[  216] = 255;
assign img[  217] = 255;
assign img[  218] = 255;
assign img[  219] = 255;
assign img[  220] = 255;
assign img[  221] = 255;
assign img[  222] = 255;
assign img[  223] = 255;
assign img[  224] = 255;
assign img[  225] = 255;
assign img[  226] = 255;
assign img[  227] = 255;
assign img[  228] = 255;
assign img[  229] = 255;
assign img[  230] = 255;
assign img[  231] = 255;
assign img[  232] = 255;
assign img[  233] = 255;
assign img[  234] = 255;
assign img[  235] = 255;
assign img[  236] = 255;
assign img[  237] = 255;
assign img[  238] = 255;
assign img[  239] = 255;
assign img[  240] = 255;
assign img[  241] = 255;
assign img[  242] = 255;
assign img[  243] = 255;
assign img[  244] = 255;
assign img[  245] = 255;
assign img[  246] = 255;
assign img[  247] = 255;
assign img[  248] = 255;
assign img[  249] = 255;
assign img[  250] = 255;
assign img[  251] = 255;
assign img[  252] = 255;
assign img[  253] = 255;
assign img[  254] = 255;
assign img[  255] = 255;
assign img[  256] = 255;
assign img[  257] = 255;
assign img[  258] = 255;
assign img[  259] = 255;
assign img[  260] = 255;
assign img[  261] = 255;
assign img[  262] = 255;
assign img[  263] = 255;
assign img[  264] = 255;
assign img[  265] = 255;
assign img[  266] = 255;
assign img[  267] = 255;
assign img[  268] = 255;
assign img[  269] = 255;
assign img[  270] = 255;
assign img[  271] = 255;
assign img[  272] = 255;
assign img[  273] = 255;
assign img[  274] = 255;
assign img[  275] = 255;
assign img[  276] = 255;
assign img[  277] = 255;
assign img[  278] = 255;
assign img[  279] = 255;
assign img[  280] = 255;
assign img[  281] = 255;
assign img[  282] = 255;
assign img[  283] = 255;
assign img[  284] = 255;
assign img[  285] = 255;
assign img[  286] = 255;
assign img[  287] = 255;
assign img[  288] = 255;
assign img[  289] = 255;
assign img[  290] = 255;
assign img[  291] = 255;
assign img[  292] = 255;
assign img[  293] = 255;
assign img[  294] = 255;
assign img[  295] = 255;
assign img[  296] = 255;
assign img[  297] = 255;
assign img[  298] = 255;
assign img[  299] = 255;
assign img[  300] = 255;
assign img[  301] = 255;
assign img[  302] = 255;
assign img[  303] = 255;
assign img[  304] = 255;
assign img[  305] = 255;
assign img[  306] = 255;
assign img[  307] = 255;
assign img[  308] = 255;
assign img[  309] = 255;
assign img[  310] = 255;
assign img[  311] = 255;
assign img[  312] = 255;
assign img[  313] = 255;
assign img[  314] = 255;
assign img[  315] = 255;
assign img[  316] = 255;
assign img[  317] = 255;
assign img[  318] = 255;
assign img[  319] = 255;
assign img[  320] = 255;
assign img[  321] = 255;
assign img[  322] = 255;
assign img[  323] = 255;
assign img[  324] = 255;
assign img[  325] = 255;
assign img[  326] = 255;
assign img[  327] = 255;
assign img[  328] = 255;
assign img[  329] = 255;
assign img[  330] = 255;
assign img[  331] = 255;
assign img[  332] = 255;
assign img[  333] = 255;
assign img[  334] = 255;
assign img[  335] = 255;
assign img[  336] = 255;
assign img[  337] = 255;
assign img[  338] = 255;
assign img[  339] = 255;
assign img[  340] = 255;
assign img[  341] = 255;
assign img[  342] = 255;
assign img[  343] = 255;
assign img[  344] = 255;
assign img[  345] = 255;
assign img[  346] = 255;
assign img[  347] = 255;
assign img[  348] = 255;
assign img[  349] = 255;
assign img[  350] = 255;
assign img[  351] = 255;
assign img[  352] = 255;
assign img[  353] = 255;
assign img[  354] = 255;
assign img[  355] = 255;
assign img[  356] = 255;
assign img[  357] = 255;
assign img[  358] = 255;
assign img[  359] = 255;
assign img[  360] = 255;
assign img[  361] = 255;
assign img[  362] = 255;
assign img[  363] = 255;
assign img[  364] = 255;
assign img[  365] = 255;
assign img[  366] = 255;
assign img[  367] = 255;
assign img[  368] = 255;
assign img[  369] = 255;
assign img[  370] = 255;
assign img[  371] = 255;
assign img[  372] = 255;
assign img[  373] = 255;
assign img[  374] = 255;
assign img[  375] = 255;
assign img[  376] = 255;
assign img[  377] = 255;
assign img[  378] = 255;
assign img[  379] = 255;
assign img[  380] = 255;
assign img[  381] = 255;
assign img[  382] = 255;
assign img[  383] = 255;
assign img[  384] = 255;
assign img[  385] = 255;
assign img[  386] = 255;
assign img[  387] = 255;
assign img[  388] = 255;
assign img[  389] = 255;
assign img[  390] = 255;
assign img[  391] = 255;
assign img[  392] = 255;
assign img[  393] = 255;
assign img[  394] = 255;
assign img[  395] = 255;
assign img[  396] = 255;
assign img[  397] = 255;
assign img[  398] = 255;
assign img[  399] = 255;
assign img[  400] = 255;
assign img[  401] = 255;
assign img[  402] = 255;
assign img[  403] = 255;
assign img[  404] = 255;
assign img[  405] = 255;
assign img[  406] = 255;
assign img[  407] = 255;
assign img[  408] = 255;
assign img[  409] = 255;
assign img[  410] = 255;
assign img[  411] = 255;
assign img[  412] = 255;
assign img[  413] = 255;
assign img[  414] = 255;
assign img[  415] = 255;
assign img[  416] = 255;
assign img[  417] = 255;
assign img[  418] = 255;
assign img[  419] = 255;
assign img[  420] = 255;
assign img[  421] = 255;
assign img[  422] = 255;
assign img[  423] = 255;
assign img[  424] = 255;
assign img[  425] = 255;
assign img[  426] = 255;
assign img[  427] = 255;
assign img[  428] = 255;
assign img[  429] = 255;
assign img[  430] = 255;
assign img[  431] = 255;
assign img[  432] = 255;
assign img[  433] = 255;
assign img[  434] = 255;
assign img[  435] = 255;
assign img[  436] = 255;
assign img[  437] = 255;
assign img[  438] = 255;
assign img[  439] = 255;
assign img[  440] = 255;
assign img[  441] = 255;
assign img[  442] = 255;
assign img[  443] = 255;
assign img[  444] = 255;
assign img[  445] = 255;
assign img[  446] = 255;
assign img[  447] = 255;
assign img[  448] = 255;
assign img[  449] = 255;
assign img[  450] = 255;
assign img[  451] = 255;
assign img[  452] = 255;
assign img[  453] = 255;
assign img[  454] = 255;
assign img[  455] = 255;
assign img[  456] = 255;
assign img[  457] = 255;
assign img[  458] = 255;
assign img[  459] = 255;
assign img[  460] = 255;
assign img[  461] = 255;
assign img[  462] = 255;
assign img[  463] = 255;
assign img[  464] = 255;
assign img[  465] = 255;
assign img[  466] = 255;
assign img[  467] = 255;
assign img[  468] = 255;
assign img[  469] = 255;
assign img[  470] = 255;
assign img[  471] = 255;
assign img[  472] = 255;
assign img[  473] = 255;
assign img[  474] = 255;
assign img[  475] = 255;
assign img[  476] = 255;
assign img[  477] = 255;
assign img[  478] = 255;
assign img[  479] = 255;
assign img[  480] = 255;
assign img[  481] = 255;
assign img[  482] = 255;
assign img[  483] = 255;
assign img[  484] = 255;
assign img[  485] = 255;
assign img[  486] = 255;
assign img[  487] = 255;
assign img[  488] = 255;
assign img[  489] = 255;
assign img[  490] = 255;
assign img[  491] = 255;
assign img[  492] = 255;
assign img[  493] = 255;
assign img[  494] = 255;
assign img[  495] = 255;
assign img[  496] = 255;
assign img[  497] = 255;
assign img[  498] = 255;
assign img[  499] = 255;
assign img[  500] = 255;
assign img[  501] = 255;
assign img[  502] = 255;
assign img[  503] = 255;
assign img[  504] = 255;
assign img[  505] = 255;
assign img[  506] = 255;
assign img[  507] = 255;
assign img[  508] = 255;
assign img[  509] = 255;
assign img[  510] = 255;
assign img[  511] = 255;
assign img[  512] = 255;
assign img[  513] = 255;
assign img[  514] = 255;
assign img[  515] = 255;
assign img[  516] = 255;
assign img[  517] = 255;
assign img[  518] = 255;
assign img[  519] = 255;
assign img[  520] = 255;
assign img[  521] = 255;
assign img[  522] = 255;
assign img[  523] = 255;
assign img[  524] = 255;
assign img[  525] = 255;
assign img[  526] = 255;
assign img[  527] = 255;
assign img[  528] = 255;
assign img[  529] = 255;
assign img[  530] = 255;
assign img[  531] = 255;
assign img[  532] = 255;
assign img[  533] = 255;
assign img[  534] = 255;
assign img[  535] = 255;
assign img[  536] = 255;
assign img[  537] = 255;
assign img[  538] = 255;
assign img[  539] = 255;
assign img[  540] = 255;
assign img[  541] = 255;
assign img[  542] = 255;
assign img[  543] = 255;
assign img[  544] = 255;
assign img[  545] = 255;
assign img[  546] = 255;
assign img[  547] = 255;
assign img[  548] = 255;
assign img[  549] = 255;
assign img[  550] = 255;
assign img[  551] = 255;
assign img[  552] = 255;
assign img[  553] = 255;
assign img[  554] = 255;
assign img[  555] = 255;
assign img[  556] = 255;
assign img[  557] = 255;
assign img[  558] = 255;
assign img[  559] = 255;
assign img[  560] = 255;
assign img[  561] = 255;
assign img[  562] = 255;
assign img[  563] = 255;
assign img[  564] = 255;
assign img[  565] = 255;
assign img[  566] = 255;
assign img[  567] = 255;
assign img[  568] = 255;
assign img[  569] = 255;
assign img[  570] = 255;
assign img[  571] = 255;
assign img[  572] = 255;
assign img[  573] = 255;
assign img[  574] = 255;
assign img[  575] = 255;
assign img[  576] = 255;
assign img[  577] = 255;
assign img[  578] = 255;
assign img[  579] = 255;
assign img[  580] = 255;
assign img[  581] = 255;
assign img[  582] = 255;
assign img[  583] = 255;
assign img[  584] = 255;
assign img[  585] = 255;
assign img[  586] = 255;
assign img[  587] = 255;
assign img[  588] = 255;
assign img[  589] = 255;
assign img[  590] = 255;
assign img[  591] = 255;
assign img[  592] = 255;
assign img[  593] = 255;
assign img[  594] = 255;
assign img[  595] = 255;
assign img[  596] = 255;
assign img[  597] = 255;
assign img[  598] = 255;
assign img[  599] = 255;
assign img[  600] = 255;
assign img[  601] = 255;
assign img[  602] = 255;
assign img[  603] = 255;
assign img[  604] = 255;
assign img[  605] = 255;
assign img[  606] = 255;
assign img[  607] = 255;
assign img[  608] = 255;
assign img[  609] = 255;
assign img[  610] = 255;
assign img[  611] = 255;
assign img[  612] = 255;
assign img[  613] = 255;
assign img[  614] = 255;
assign img[  615] = 255;
assign img[  616] = 255;
assign img[  617] = 255;
assign img[  618] = 255;
assign img[  619] = 255;
assign img[  620] = 255;
assign img[  621] = 255;
assign img[  622] = 255;
assign img[  623] = 255;
assign img[  624] = 255;
assign img[  625] = 255;
assign img[  626] = 255;
assign img[  627] = 255;
assign img[  628] = 255;
assign img[  629] = 255;
assign img[  630] = 255;
assign img[  631] = 255;
assign img[  632] = 255;
assign img[  633] = 255;
assign img[  634] = 255;
assign img[  635] = 255;
assign img[  636] = 255;
assign img[  637] = 255;
assign img[  638] = 255;
assign img[  639] = 255;
assign img[  640] = 255;
assign img[  641] = 255;
assign img[  642] = 255;
assign img[  643] = 255;
assign img[  644] = 255;
assign img[  645] = 255;
assign img[  646] = 255;
assign img[  647] = 255;
assign img[  648] = 255;
assign img[  649] = 255;
assign img[  650] = 255;
assign img[  651] = 255;
assign img[  652] = 255;
assign img[  653] = 255;
assign img[  654] = 255;
assign img[  655] = 255;
assign img[  656] = 255;
assign img[  657] = 255;
assign img[  658] = 255;
assign img[  659] = 255;
assign img[  660] = 255;
assign img[  661] = 255;
assign img[  662] = 255;
assign img[  663] = 255;
assign img[  664] = 255;
assign img[  665] = 255;
assign img[  666] = 255;
assign img[  667] = 255;
assign img[  668] = 255;
assign img[  669] = 255;
assign img[  670] = 255;
assign img[  671] = 255;
assign img[  672] = 255;
assign img[  673] = 255;
assign img[  674] = 255;
assign img[  675] = 255;
assign img[  676] = 255;
assign img[  677] = 255;
assign img[  678] = 255;
assign img[  679] = 255;
assign img[  680] = 255;
assign img[  681] = 255;
assign img[  682] = 255;
assign img[  683] = 255;
assign img[  684] = 255;
assign img[  685] = 255;
assign img[  686] = 255;
assign img[  687] = 255;
assign img[  688] = 255;
assign img[  689] = 255;
assign img[  690] = 255;
assign img[  691] = 255;
assign img[  692] = 255;
assign img[  693] = 255;
assign img[  694] = 255;
assign img[  695] = 255;
assign img[  696] = 255;
assign img[  697] = 255;
assign img[  698] = 255;
assign img[  699] = 255;
assign img[  700] = 255;
assign img[  701] = 255;
assign img[  702] = 255;
assign img[  703] = 255;
assign img[  704] = 255;
assign img[  705] = 255;
assign img[  706] = 255;
assign img[  707] = 255;
assign img[  708] = 255;
assign img[  709] = 255;
assign img[  710] = 255;
assign img[  711] = 255;
assign img[  712] = 255;
assign img[  713] = 255;
assign img[  714] = 255;
assign img[  715] = 255;
assign img[  716] = 255;
assign img[  717] = 255;
assign img[  718] = 255;
assign img[  719] = 255;
assign img[  720] = 255;
assign img[  721] = 255;
assign img[  722] = 255;
assign img[  723] = 255;
assign img[  724] = 255;
assign img[  725] = 255;
assign img[  726] = 255;
assign img[  727] = 255;
assign img[  728] = 255;
assign img[  729] = 255;
assign img[  730] = 255;
assign img[  731] = 255;
assign img[  732] = 255;
assign img[  733] = 255;
assign img[  734] = 255;
assign img[  735] = 255;
assign img[  736] = 255;
assign img[  737] = 255;
assign img[  738] = 255;
assign img[  739] = 255;
assign img[  740] = 255;
assign img[  741] = 255;
assign img[  742] = 255;
assign img[  743] = 255;
assign img[  744] = 255;
assign img[  745] = 255;
assign img[  746] = 255;
assign img[  747] = 255;
assign img[  748] = 255;
assign img[  749] = 255;
assign img[  750] = 255;
assign img[  751] = 255;
assign img[  752] = 255;
assign img[  753] = 255;
assign img[  754] = 255;
assign img[  755] = 255;
assign img[  756] = 255;
assign img[  757] = 255;
assign img[  758] = 255;
assign img[  759] = 255;
assign img[  760] = 255;
assign img[  761] = 255;
assign img[  762] = 255;
assign img[  763] = 255;
assign img[  764] = 255;
assign img[  765] = 255;
assign img[  766] = 255;
assign img[  767] = 255;
assign img[  768] = 255;
assign img[  769] = 255;
assign img[  770] = 255;
assign img[  771] = 255;
assign img[  772] = 255;
assign img[  773] = 255;
assign img[  774] = 255;
assign img[  775] = 255;
assign img[  776] = 255;
assign img[  777] = 255;
assign img[  778] = 255;
assign img[  779] = 255;
assign img[  780] = 255;
assign img[  781] = 255;
assign img[  782] = 255;
assign img[  783] = 255;
assign img[  784] = 255;
assign img[  785] = 255;
assign img[  786] = 255;
assign img[  787] = 255;
assign img[  788] = 255;
assign img[  789] = 255;
assign img[  790] = 255;
assign img[  791] = 255;
assign img[  792] = 255;
assign img[  793] = 255;
assign img[  794] = 255;
assign img[  795] = 255;
assign img[  796] = 255;
assign img[  797] = 255;
assign img[  798] = 255;
assign img[  799] = 255;
assign img[  800] = 255;
assign img[  801] = 255;
assign img[  802] = 255;
assign img[  803] = 255;
assign img[  804] = 255;
assign img[  805] = 255;
assign img[  806] = 255;
assign img[  807] = 255;
assign img[  808] = 255;
assign img[  809] = 255;
assign img[  810] = 255;
assign img[  811] = 255;
assign img[  812] = 255;
assign img[  813] = 255;
assign img[  814] = 255;
assign img[  815] = 255;
assign img[  816] = 255;
assign img[  817] = 255;
assign img[  818] = 255;
assign img[  819] = 255;
assign img[  820] = 255;
assign img[  821] = 255;
assign img[  822] = 255;
assign img[  823] = 255;
assign img[  824] = 255;
assign img[  825] = 255;
assign img[  826] = 255;
assign img[  827] = 255;
assign img[  828] = 255;
assign img[  829] = 255;
assign img[  830] = 255;
assign img[  831] = 255;
assign img[  832] = 255;
assign img[  833] = 255;
assign img[  834] = 255;
assign img[  835] = 255;
assign img[  836] = 255;
assign img[  837] = 255;
assign img[  838] = 255;
assign img[  839] = 255;
assign img[  840] = 255;
assign img[  841] = 255;
assign img[  842] = 255;
assign img[  843] = 255;
assign img[  844] = 255;
assign img[  845] = 255;
assign img[  846] = 255;
assign img[  847] = 255;
assign img[  848] = 255;
assign img[  849] = 255;
assign img[  850] = 255;
assign img[  851] = 255;
assign img[  852] = 255;
assign img[  853] = 255;
assign img[  854] = 255;
assign img[  855] = 255;
assign img[  856] = 255;
assign img[  857] = 255;
assign img[  858] = 255;
assign img[  859] = 255;
assign img[  860] = 255;
assign img[  861] = 255;
assign img[  862] = 255;
assign img[  863] = 255;
assign img[  864] = 255;
assign img[  865] = 255;
assign img[  866] = 255;
assign img[  867] = 255;
assign img[  868] = 255;
assign img[  869] = 255;
assign img[  870] = 255;
assign img[  871] = 255;
assign img[  872] = 255;
assign img[  873] = 255;
assign img[  874] = 255;
assign img[  875] = 255;
assign img[  876] = 255;
assign img[  877] = 255;
assign img[  878] = 255;
assign img[  879] = 255;
assign img[  880] = 255;
assign img[  881] = 255;
assign img[  882] = 255;
assign img[  883] = 255;
assign img[  884] = 255;
assign img[  885] = 255;
assign img[  886] = 255;
assign img[  887] = 255;
assign img[  888] = 255;
assign img[  889] = 255;
assign img[  890] = 255;
assign img[  891] = 255;
assign img[  892] = 255;
assign img[  893] = 255;
assign img[  894] = 255;
assign img[  895] = 255;
assign img[  896] = 255;
assign img[  897] = 255;
assign img[  898] = 255;
assign img[  899] = 255;
assign img[  900] = 255;
assign img[  901] = 255;
assign img[  902] = 255;
assign img[  903] = 255;
assign img[  904] = 255;
assign img[  905] = 255;
assign img[  906] = 255;
assign img[  907] = 255;
assign img[  908] = 255;
assign img[  909] = 255;
assign img[  910] = 255;
assign img[  911] = 255;
assign img[  912] = 255;
assign img[  913] = 255;
assign img[  914] = 255;
assign img[  915] = 255;
assign img[  916] = 255;
assign img[  917] = 255;
assign img[  918] = 255;
assign img[  919] = 255;
assign img[  920] = 255;
assign img[  921] = 255;
assign img[  922] = 255;
assign img[  923] = 255;
assign img[  924] = 255;
assign img[  925] = 255;
assign img[  926] = 255;
assign img[  927] = 255;
assign img[  928] = 255;
assign img[  929] = 255;
assign img[  930] = 255;
assign img[  931] = 255;
assign img[  932] = 255;
assign img[  933] = 255;
assign img[  934] = 255;
assign img[  935] = 255;
assign img[  936] = 255;
assign img[  937] = 255;
assign img[  938] = 255;
assign img[  939] = 255;
assign img[  940] = 255;
assign img[  941] = 255;
assign img[  942] = 255;
assign img[  943] = 255;
assign img[  944] = 255;
assign img[  945] = 255;
assign img[  946] = 255;
assign img[  947] = 255;
assign img[  948] = 255;
assign img[  949] = 255;
assign img[  950] = 255;
assign img[  951] = 255;
assign img[  952] = 255;
assign img[  953] = 255;
assign img[  954] = 255;
assign img[  955] = 255;
assign img[  956] = 255;
assign img[  957] = 255;
assign img[  958] = 255;
assign img[  959] = 255;
assign img[  960] = 255;
assign img[  961] = 255;
assign img[  962] = 255;
assign img[  963] = 255;
assign img[  964] = 255;
assign img[  965] = 255;
assign img[  966] = 255;
assign img[  967] = 255;
assign img[  968] = 255;
assign img[  969] = 255;
assign img[  970] = 255;
assign img[  971] = 255;
assign img[  972] = 255;
assign img[  973] = 255;
assign img[  974] = 255;
assign img[  975] = 255;
assign img[  976] = 255;
assign img[  977] = 255;
assign img[  978] = 255;
assign img[  979] = 255;
assign img[  980] = 255;
assign img[  981] = 255;
assign img[  982] = 255;
assign img[  983] = 255;
assign img[  984] = 255;
assign img[  985] = 255;
assign img[  986] = 255;
assign img[  987] = 255;
assign img[  988] = 255;
assign img[  989] = 255;
assign img[  990] = 255;
assign img[  991] = 255;
assign img[  992] = 255;
assign img[  993] = 255;
assign img[  994] = 255;
assign img[  995] = 255;
assign img[  996] = 255;
assign img[  997] = 255;
assign img[  998] = 255;
assign img[  999] = 255;
assign img[ 1000] = 255;
assign img[ 1001] = 255;
assign img[ 1002] = 255;
assign img[ 1003] = 255;
assign img[ 1004] = 255;
assign img[ 1005] = 255;
assign img[ 1006] = 255;
assign img[ 1007] = 255;
assign img[ 1008] = 255;
assign img[ 1009] = 255;
assign img[ 1010] = 255;
assign img[ 1011] = 255;
assign img[ 1012] = 255;
assign img[ 1013] = 255;
assign img[ 1014] = 255;
assign img[ 1015] = 255;
assign img[ 1016] = 255;
assign img[ 1017] = 255;
assign img[ 1018] = 255;
assign img[ 1019] = 255;
assign img[ 1020] = 255;
assign img[ 1021] = 255;
assign img[ 1022] = 255;
assign img[ 1023] = 255;
assign img[ 1024] = 255;
assign img[ 1025] = 255;
assign img[ 1026] = 255;
assign img[ 1027] = 255;
assign img[ 1028] = 255;
assign img[ 1029] = 255;
assign img[ 1030] = 255;
assign img[ 1031] = 255;
assign img[ 1032] = 255;
assign img[ 1033] = 255;
assign img[ 1034] = 255;
assign img[ 1035] = 255;
assign img[ 1036] = 255;
assign img[ 1037] = 255;
assign img[ 1038] = 255;
assign img[ 1039] = 255;
assign img[ 1040] = 255;
assign img[ 1041] = 255;
assign img[ 1042] = 255;
assign img[ 1043] = 255;
assign img[ 1044] = 255;
assign img[ 1045] = 255;
assign img[ 1046] = 255;
assign img[ 1047] = 255;
assign img[ 1048] = 255;
assign img[ 1049] = 255;
assign img[ 1050] = 255;
assign img[ 1051] = 255;
assign img[ 1052] = 255;
assign img[ 1053] = 255;
assign img[ 1054] = 255;
assign img[ 1055] = 255;
assign img[ 1056] = 255;
assign img[ 1057] = 255;
assign img[ 1058] = 255;
assign img[ 1059] = 255;
assign img[ 1060] = 255;
assign img[ 1061] = 255;
assign img[ 1062] = 255;
assign img[ 1063] = 255;
assign img[ 1064] = 255;
assign img[ 1065] = 255;
assign img[ 1066] = 255;
assign img[ 1067] = 255;
assign img[ 1068] = 255;
assign img[ 1069] = 255;
assign img[ 1070] = 255;
assign img[ 1071] = 255;
assign img[ 1072] = 255;
assign img[ 1073] = 255;
assign img[ 1074] = 255;
assign img[ 1075] = 255;
assign img[ 1076] = 255;
assign img[ 1077] = 255;
assign img[ 1078] = 255;
assign img[ 1079] = 255;
assign img[ 1080] = 255;
assign img[ 1081] = 255;
assign img[ 1082] = 255;
assign img[ 1083] = 255;
assign img[ 1084] = 255;
assign img[ 1085] = 255;
assign img[ 1086] = 255;
assign img[ 1087] = 255;
assign img[ 1088] = 255;
assign img[ 1089] = 255;
assign img[ 1090] = 255;
assign img[ 1091] = 255;
assign img[ 1092] = 255;
assign img[ 1093] = 255;
assign img[ 1094] = 255;
assign img[ 1095] = 255;
assign img[ 1096] = 255;
assign img[ 1097] = 255;
assign img[ 1098] = 255;
assign img[ 1099] = 255;
assign img[ 1100] = 255;
assign img[ 1101] = 255;
assign img[ 1102] = 255;
assign img[ 1103] = 255;
assign img[ 1104] = 255;
assign img[ 1105] = 255;
assign img[ 1106] = 255;
assign img[ 1107] = 255;
assign img[ 1108] = 255;
assign img[ 1109] = 255;
assign img[ 1110] = 255;
assign img[ 1111] = 255;
assign img[ 1112] = 255;
assign img[ 1113] = 255;
assign img[ 1114] = 255;
assign img[ 1115] = 255;
assign img[ 1116] = 255;
assign img[ 1117] = 255;
assign img[ 1118] = 255;
assign img[ 1119] = 255;
assign img[ 1120] = 255;
assign img[ 1121] = 255;
assign img[ 1122] = 255;
assign img[ 1123] = 255;
assign img[ 1124] = 255;
assign img[ 1125] = 255;
assign img[ 1126] = 255;
assign img[ 1127] = 255;
assign img[ 1128] = 255;
assign img[ 1129] = 255;
assign img[ 1130] = 255;
assign img[ 1131] = 255;
assign img[ 1132] = 255;
assign img[ 1133] = 255;
assign img[ 1134] = 255;
assign img[ 1135] = 255;
assign img[ 1136] = 255;
assign img[ 1137] = 255;
assign img[ 1138] = 255;
assign img[ 1139] = 255;
assign img[ 1140] = 255;
assign img[ 1141] = 255;
assign img[ 1142] = 255;
assign img[ 1143] = 255;
assign img[ 1144] = 255;
assign img[ 1145] = 255;
assign img[ 1146] = 255;
assign img[ 1147] = 255;
assign img[ 1148] = 255;
assign img[ 1149] = 255;
assign img[ 1150] = 255;
assign img[ 1151] = 255;
assign img[ 1152] = 255;
assign img[ 1153] = 255;
assign img[ 1154] = 255;
assign img[ 1155] = 255;
assign img[ 1156] = 255;
assign img[ 1157] = 255;
assign img[ 1158] = 255;
assign img[ 1159] = 255;
assign img[ 1160] = 255;
assign img[ 1161] = 255;
assign img[ 1162] = 255;
assign img[ 1163] = 255;
assign img[ 1164] = 255;
assign img[ 1165] = 255;
assign img[ 1166] = 255;
assign img[ 1167] = 255;
assign img[ 1168] = 255;
assign img[ 1169] = 255;
assign img[ 1170] = 255;
assign img[ 1171] = 255;
assign img[ 1172] = 255;
assign img[ 1173] = 255;
assign img[ 1174] = 255;
assign img[ 1175] = 255;
assign img[ 1176] = 255;
assign img[ 1177] = 255;
assign img[ 1178] = 255;
assign img[ 1179] = 255;
assign img[ 1180] = 255;
assign img[ 1181] = 255;
assign img[ 1182] = 255;
assign img[ 1183] = 255;
assign img[ 1184] = 255;
assign img[ 1185] = 255;
assign img[ 1186] = 255;
assign img[ 1187] = 255;
assign img[ 1188] = 255;
assign img[ 1189] = 255;
assign img[ 1190] = 255;
assign img[ 1191] = 255;
assign img[ 1192] = 255;
assign img[ 1193] = 255;
assign img[ 1194] = 255;
assign img[ 1195] = 255;
assign img[ 1196] = 255;
assign img[ 1197] = 255;
assign img[ 1198] = 255;
assign img[ 1199] = 255;
assign img[ 1200] = 255;
assign img[ 1201] = 255;
assign img[ 1202] = 255;
assign img[ 1203] = 255;
assign img[ 1204] = 255;
assign img[ 1205] = 255;
assign img[ 1206] = 255;
assign img[ 1207] = 255;
assign img[ 1208] = 255;
assign img[ 1209] = 255;
assign img[ 1210] = 255;
assign img[ 1211] = 255;
assign img[ 1212] = 255;
assign img[ 1213] = 255;
assign img[ 1214] = 255;
assign img[ 1215] = 255;
assign img[ 1216] = 255;
assign img[ 1217] = 255;
assign img[ 1218] = 255;
assign img[ 1219] = 255;
assign img[ 1220] = 255;
assign img[ 1221] = 255;
assign img[ 1222] = 255;
assign img[ 1223] = 255;
assign img[ 1224] = 255;
assign img[ 1225] = 255;
assign img[ 1226] = 255;
assign img[ 1227] = 255;
assign img[ 1228] = 255;
assign img[ 1229] = 255;
assign img[ 1230] = 255;
assign img[ 1231] = 255;
assign img[ 1232] = 255;
assign img[ 1233] = 255;
assign img[ 1234] = 255;
assign img[ 1235] = 255;
assign img[ 1236] = 255;
assign img[ 1237] = 255;
assign img[ 1238] = 255;
assign img[ 1239] = 255;
assign img[ 1240] = 255;
assign img[ 1241] = 255;
assign img[ 1242] = 255;
assign img[ 1243] = 255;
assign img[ 1244] = 255;
assign img[ 1245] = 255;
assign img[ 1246] = 255;
assign img[ 1247] = 255;
assign img[ 1248] = 255;
assign img[ 1249] = 255;
assign img[ 1250] = 255;
assign img[ 1251] = 255;
assign img[ 1252] = 255;
assign img[ 1253] = 255;
assign img[ 1254] = 255;
assign img[ 1255] = 255;
assign img[ 1256] = 255;
assign img[ 1257] = 255;
assign img[ 1258] = 255;
assign img[ 1259] = 255;
assign img[ 1260] = 255;
assign img[ 1261] = 255;
assign img[ 1262] = 255;
assign img[ 1263] = 255;
assign img[ 1264] = 255;
assign img[ 1265] = 255;
assign img[ 1266] = 255;
assign img[ 1267] = 255;
assign img[ 1268] = 255;
assign img[ 1269] = 255;
assign img[ 1270] = 255;
assign img[ 1271] = 255;
assign img[ 1272] = 255;
assign img[ 1273] = 255;
assign img[ 1274] = 255;
assign img[ 1275] = 255;
assign img[ 1276] = 255;
assign img[ 1277] = 255;
assign img[ 1278] = 255;
assign img[ 1279] = 255;
assign img[ 1280] = 255;
assign img[ 1281] = 255;
assign img[ 1282] = 255;
assign img[ 1283] = 255;
assign img[ 1284] = 255;
assign img[ 1285] = 255;
assign img[ 1286] = 255;
assign img[ 1287] = 255;
assign img[ 1288] = 255;
assign img[ 1289] = 255;
assign img[ 1290] = 255;
assign img[ 1291] = 255;
assign img[ 1292] = 255;
assign img[ 1293] = 255;
assign img[ 1294] = 255;
assign img[ 1295] = 255;
assign img[ 1296] = 255;
assign img[ 1297] = 255;
assign img[ 1298] = 255;
assign img[ 1299] = 255;
assign img[ 1300] = 255;
assign img[ 1301] = 255;
assign img[ 1302] = 255;
assign img[ 1303] = 255;
assign img[ 1304] = 255;
assign img[ 1305] = 255;
assign img[ 1306] = 255;
assign img[ 1307] = 255;
assign img[ 1308] = 255;
assign img[ 1309] = 255;
assign img[ 1310] = 255;
assign img[ 1311] = 255;
assign img[ 1312] = 255;
assign img[ 1313] = 255;
assign img[ 1314] = 255;
assign img[ 1315] = 255;
assign img[ 1316] = 255;
assign img[ 1317] = 255;
assign img[ 1318] = 255;
assign img[ 1319] = 255;
assign img[ 1320] = 255;
assign img[ 1321] = 255;
assign img[ 1322] = 255;
assign img[ 1323] = 255;
assign img[ 1324] = 255;
assign img[ 1325] = 255;
assign img[ 1326] = 255;
assign img[ 1327] = 255;
assign img[ 1328] = 255;
assign img[ 1329] = 255;
assign img[ 1330] = 255;
assign img[ 1331] = 255;
assign img[ 1332] = 255;
assign img[ 1333] = 255;
assign img[ 1334] = 255;
assign img[ 1335] = 255;
assign img[ 1336] = 255;
assign img[ 1337] = 255;
assign img[ 1338] = 255;
assign img[ 1339] = 255;
assign img[ 1340] = 255;
assign img[ 1341] = 255;
assign img[ 1342] = 255;
assign img[ 1343] = 255;
assign img[ 1344] = 255;
assign img[ 1345] = 255;
assign img[ 1346] = 255;
assign img[ 1347] = 255;
assign img[ 1348] = 255;
assign img[ 1349] = 255;
assign img[ 1350] = 255;
assign img[ 1351] = 255;
assign img[ 1352] = 255;
assign img[ 1353] = 255;
assign img[ 1354] = 255;
assign img[ 1355] = 255;
assign img[ 1356] = 255;
assign img[ 1357] = 255;
assign img[ 1358] = 255;
assign img[ 1359] = 255;
assign img[ 1360] = 255;
assign img[ 1361] = 255;
assign img[ 1362] = 255;
assign img[ 1363] = 255;
assign img[ 1364] = 255;
assign img[ 1365] = 255;
assign img[ 1366] = 255;
assign img[ 1367] = 255;
assign img[ 1368] = 255;
assign img[ 1369] = 255;
assign img[ 1370] = 255;
assign img[ 1371] = 255;
assign img[ 1372] = 255;
assign img[ 1373] = 255;
assign img[ 1374] = 255;
assign img[ 1375] = 255;
assign img[ 1376] = 255;
assign img[ 1377] = 255;
assign img[ 1378] = 255;
assign img[ 1379] = 255;
assign img[ 1380] = 255;
assign img[ 1381] = 255;
assign img[ 1382] = 255;
assign img[ 1383] = 255;
assign img[ 1384] = 255;
assign img[ 1385] = 255;
assign img[ 1386] = 255;
assign img[ 1387] = 255;
assign img[ 1388] = 255;
assign img[ 1389] = 255;
assign img[ 1390] = 255;
assign img[ 1391] = 255;
assign img[ 1392] = 255;
assign img[ 1393] = 255;
assign img[ 1394] = 255;
assign img[ 1395] = 255;
assign img[ 1396] = 255;
assign img[ 1397] = 255;
assign img[ 1398] = 255;
assign img[ 1399] = 255;
assign img[ 1400] = 255;
assign img[ 1401] = 255;
assign img[ 1402] = 255;
assign img[ 1403] = 255;
assign img[ 1404] = 255;
assign img[ 1405] = 255;
assign img[ 1406] = 255;
assign img[ 1407] = 255;
assign img[ 1408] = 255;
assign img[ 1409] = 255;
assign img[ 1410] = 255;
assign img[ 1411] = 255;
assign img[ 1412] = 255;
assign img[ 1413] = 255;
assign img[ 1414] = 255;
assign img[ 1415] = 255;
assign img[ 1416] = 255;
assign img[ 1417] = 255;
assign img[ 1418] = 255;
assign img[ 1419] = 255;
assign img[ 1420] = 255;
assign img[ 1421] = 255;
assign img[ 1422] = 255;
assign img[ 1423] = 255;
assign img[ 1424] = 255;
assign img[ 1425] = 255;
assign img[ 1426] = 255;
assign img[ 1427] = 255;
assign img[ 1428] = 255;
assign img[ 1429] = 255;
assign img[ 1430] = 255;
assign img[ 1431] = 255;
assign img[ 1432] = 255;
assign img[ 1433] = 255;
assign img[ 1434] = 255;
assign img[ 1435] = 255;
assign img[ 1436] = 255;
assign img[ 1437] = 255;
assign img[ 1438] = 255;
assign img[ 1439] = 255;
assign img[ 1440] = 255;
assign img[ 1441] = 255;
assign img[ 1442] = 255;
assign img[ 1443] = 255;
assign img[ 1444] = 255;
assign img[ 1445] = 255;
assign img[ 1446] = 255;
assign img[ 1447] = 255;
assign img[ 1448] = 255;
assign img[ 1449] = 255;
assign img[ 1450] = 255;
assign img[ 1451] = 255;
assign img[ 1452] = 255;
assign img[ 1453] = 255;
assign img[ 1454] = 255;
assign img[ 1455] = 255;
assign img[ 1456] = 255;
assign img[ 1457] = 255;
assign img[ 1458] = 255;
assign img[ 1459] = 255;
assign img[ 1460] = 255;
assign img[ 1461] = 255;
assign img[ 1462] = 255;
assign img[ 1463] = 255;
assign img[ 1464] = 255;
assign img[ 1465] = 255;
assign img[ 1466] = 255;
assign img[ 1467] = 255;
assign img[ 1468] = 255;
assign img[ 1469] = 255;
assign img[ 1470] = 255;
assign img[ 1471] = 255;
assign img[ 1472] = 255;
assign img[ 1473] = 255;
assign img[ 1474] = 255;
assign img[ 1475] = 255;
assign img[ 1476] = 255;
assign img[ 1477] = 255;
assign img[ 1478] = 255;
assign img[ 1479] = 255;
assign img[ 1480] = 255;
assign img[ 1481] = 255;
assign img[ 1482] = 255;
assign img[ 1483] = 255;
assign img[ 1484] = 255;
assign img[ 1485] = 255;
assign img[ 1486] = 255;
assign img[ 1487] = 255;
assign img[ 1488] = 255;
assign img[ 1489] = 255;
assign img[ 1490] = 255;
assign img[ 1491] = 255;
assign img[ 1492] = 255;
assign img[ 1493] = 255;
assign img[ 1494] = 255;
assign img[ 1495] = 255;
assign img[ 1496] = 255;
assign img[ 1497] = 255;
assign img[ 1498] = 255;
assign img[ 1499] = 255;
assign img[ 1500] = 255;
assign img[ 1501] = 255;
assign img[ 1502] = 255;
assign img[ 1503] = 255;
assign img[ 1504] = 255;
assign img[ 1505] = 255;
assign img[ 1506] = 255;
assign img[ 1507] = 255;
assign img[ 1508] = 255;
assign img[ 1509] = 255;
assign img[ 1510] = 255;
assign img[ 1511] = 255;
assign img[ 1512] = 255;
assign img[ 1513] = 255;
assign img[ 1514] = 255;
assign img[ 1515] = 255;
assign img[ 1516] = 255;
assign img[ 1517] = 255;
assign img[ 1518] = 255;
assign img[ 1519] = 255;
assign img[ 1520] = 255;
assign img[ 1521] = 255;
assign img[ 1522] = 255;
assign img[ 1523] = 255;
assign img[ 1524] = 255;
assign img[ 1525] = 255;
assign img[ 1526] = 255;
assign img[ 1527] = 255;
assign img[ 1528] = 255;
assign img[ 1529] = 255;
assign img[ 1530] = 255;
assign img[ 1531] = 255;
assign img[ 1532] = 255;
assign img[ 1533] = 255;
assign img[ 1534] = 255;
assign img[ 1535] = 255;
assign img[ 1536] = 255;
assign img[ 1537] = 255;
assign img[ 1538] = 255;
assign img[ 1539] = 255;
assign img[ 1540] = 255;
assign img[ 1541] = 255;
assign img[ 1542] = 255;
assign img[ 1543] = 255;
assign img[ 1544] = 255;
assign img[ 1545] = 255;
assign img[ 1546] = 255;
assign img[ 1547] = 255;
assign img[ 1548] = 255;
assign img[ 1549] = 255;
assign img[ 1550] = 255;
assign img[ 1551] = 255;
assign img[ 1552] = 255;
assign img[ 1553] = 255;
assign img[ 1554] = 255;
assign img[ 1555] = 255;
assign img[ 1556] = 255;
assign img[ 1557] = 255;
assign img[ 1558] = 255;
assign img[ 1559] = 255;
assign img[ 1560] = 255;
assign img[ 1561] = 255;
assign img[ 1562] = 255;
assign img[ 1563] = 255;
assign img[ 1564] = 255;
assign img[ 1565] = 255;
assign img[ 1566] = 255;
assign img[ 1567] = 255;
assign img[ 1568] = 255;
assign img[ 1569] = 255;
assign img[ 1570] = 255;
assign img[ 1571] = 255;
assign img[ 1572] = 255;
assign img[ 1573] = 255;
assign img[ 1574] = 255;
assign img[ 1575] = 255;
assign img[ 1576] = 255;
assign img[ 1577] = 255;
assign img[ 1578] = 255;
assign img[ 1579] = 255;
assign img[ 1580] = 255;
assign img[ 1581] = 255;
assign img[ 1582] = 255;
assign img[ 1583] = 255;
assign img[ 1584] = 255;
assign img[ 1585] = 255;
assign img[ 1586] = 255;
assign img[ 1587] = 255;
assign img[ 1588] = 255;
assign img[ 1589] = 255;
assign img[ 1590] = 255;
assign img[ 1591] = 255;
assign img[ 1592] = 255;
assign img[ 1593] = 255;
assign img[ 1594] = 255;
assign img[ 1595] = 255;
assign img[ 1596] = 255;
assign img[ 1597] = 255;
assign img[ 1598] = 255;
assign img[ 1599] = 255;
assign img[ 1600] = 255;
assign img[ 1601] = 255;
assign img[ 1602] = 255;
assign img[ 1603] = 255;
assign img[ 1604] = 255;
assign img[ 1605] = 255;
assign img[ 1606] = 255;
assign img[ 1607] = 255;
assign img[ 1608] = 255;
assign img[ 1609] = 255;
assign img[ 1610] = 255;
assign img[ 1611] = 255;
assign img[ 1612] = 255;
assign img[ 1613] = 255;
assign img[ 1614] = 255;
assign img[ 1615] = 255;
assign img[ 1616] = 255;
assign img[ 1617] = 255;
assign img[ 1618] = 255;
assign img[ 1619] = 255;
assign img[ 1620] = 255;
assign img[ 1621] = 255;
assign img[ 1622] = 255;
assign img[ 1623] = 255;
assign img[ 1624] = 255;
assign img[ 1625] = 255;
assign img[ 1626] = 255;
assign img[ 1627] = 255;
assign img[ 1628] = 255;
assign img[ 1629] = 255;
assign img[ 1630] = 255;
assign img[ 1631] = 255;
assign img[ 1632] = 255;
assign img[ 1633] = 255;
assign img[ 1634] = 255;
assign img[ 1635] = 255;
assign img[ 1636] = 255;
assign img[ 1637] = 255;
assign img[ 1638] = 255;
assign img[ 1639] = 255;
assign img[ 1640] = 255;
assign img[ 1641] = 255;
assign img[ 1642] = 255;
assign img[ 1643] = 255;
assign img[ 1644] = 255;
assign img[ 1645] = 255;
assign img[ 1646] = 255;
assign img[ 1647] = 255;
assign img[ 1648] = 255;
assign img[ 1649] = 255;
assign img[ 1650] = 255;
assign img[ 1651] = 255;
assign img[ 1652] = 255;
assign img[ 1653] = 255;
assign img[ 1654] = 255;
assign img[ 1655] = 255;
assign img[ 1656] = 255;
assign img[ 1657] = 255;
assign img[ 1658] = 255;
assign img[ 1659] = 255;
assign img[ 1660] = 255;
assign img[ 1661] = 255;
assign img[ 1662] = 255;
assign img[ 1663] = 255;
assign img[ 1664] = 255;
assign img[ 1665] = 255;
assign img[ 1666] = 255;
assign img[ 1667] = 255;
assign img[ 1668] = 255;
assign img[ 1669] = 255;
assign img[ 1670] = 255;
assign img[ 1671] = 255;
assign img[ 1672] = 255;
assign img[ 1673] = 255;
assign img[ 1674] = 255;
assign img[ 1675] = 255;
assign img[ 1676] = 255;
assign img[ 1677] = 255;
assign img[ 1678] = 255;
assign img[ 1679] = 255;
assign img[ 1680] = 255;
assign img[ 1681] = 255;
assign img[ 1682] = 255;
assign img[ 1683] = 255;
assign img[ 1684] = 255;
assign img[ 1685] = 255;
assign img[ 1686] = 255;
assign img[ 1687] = 255;
assign img[ 1688] = 255;
assign img[ 1689] = 255;
assign img[ 1690] = 255;
assign img[ 1691] = 255;
assign img[ 1692] = 255;
assign img[ 1693] = 255;
assign img[ 1694] = 255;
assign img[ 1695] = 255;
assign img[ 1696] = 255;
assign img[ 1697] = 255;
assign img[ 1698] = 255;
assign img[ 1699] = 255;
assign img[ 1700] = 255;
assign img[ 1701] = 255;
assign img[ 1702] = 255;
assign img[ 1703] = 255;
assign img[ 1704] = 255;
assign img[ 1705] = 255;
assign img[ 1706] = 255;
assign img[ 1707] = 255;
assign img[ 1708] = 255;
assign img[ 1709] = 255;
assign img[ 1710] = 255;
assign img[ 1711] = 255;
assign img[ 1712] = 255;
assign img[ 1713] = 255;
assign img[ 1714] = 255;
assign img[ 1715] = 255;
assign img[ 1716] = 255;
assign img[ 1717] = 255;
assign img[ 1718] = 255;
assign img[ 1719] = 255;
assign img[ 1720] = 255;
assign img[ 1721] = 255;
assign img[ 1722] = 255;
assign img[ 1723] = 255;
assign img[ 1724] = 255;
assign img[ 1725] = 255;
assign img[ 1726] = 255;
assign img[ 1727] = 255;
assign img[ 1728] = 255;
assign img[ 1729] = 255;
assign img[ 1730] = 255;
assign img[ 1731] = 255;
assign img[ 1732] = 255;
assign img[ 1733] = 255;
assign img[ 1734] = 255;
assign img[ 1735] = 255;
assign img[ 1736] = 255;
assign img[ 1737] = 255;
assign img[ 1738] = 255;
assign img[ 1739] = 255;
assign img[ 1740] = 255;
assign img[ 1741] = 255;
assign img[ 1742] = 255;
assign img[ 1743] = 255;
assign img[ 1744] = 255;
assign img[ 1745] = 255;
assign img[ 1746] = 255;
assign img[ 1747] = 255;
assign img[ 1748] = 255;
assign img[ 1749] = 255;
assign img[ 1750] = 255;
assign img[ 1751] = 255;
assign img[ 1752] = 255;
assign img[ 1753] = 255;
assign img[ 1754] = 255;
assign img[ 1755] = 255;
assign img[ 1756] = 255;
assign img[ 1757] = 255;
assign img[ 1758] = 255;
assign img[ 1759] = 255;
assign img[ 1760] = 255;
assign img[ 1761] = 255;
assign img[ 1762] = 255;
assign img[ 1763] = 255;
assign img[ 1764] = 255;
assign img[ 1765] = 255;
assign img[ 1766] = 255;
assign img[ 1767] = 255;
assign img[ 1768] = 255;
assign img[ 1769] = 255;
assign img[ 1770] = 255;
assign img[ 1771] = 255;
assign img[ 1772] = 255;
assign img[ 1773] = 255;
assign img[ 1774] = 255;
assign img[ 1775] = 255;
assign img[ 1776] = 255;
assign img[ 1777] = 255;
assign img[ 1778] = 255;
assign img[ 1779] = 255;
assign img[ 1780] = 255;
assign img[ 1781] = 255;
assign img[ 1782] = 255;
assign img[ 1783] = 255;
assign img[ 1784] = 255;
assign img[ 1785] = 255;
assign img[ 1786] = 255;
assign img[ 1787] = 255;
assign img[ 1788] = 255;
assign img[ 1789] = 255;
assign img[ 1790] = 255;
assign img[ 1791] = 255;
assign img[ 1792] = 255;
assign img[ 1793] = 255;
assign img[ 1794] = 255;
assign img[ 1795] = 255;
assign img[ 1796] = 255;
assign img[ 1797] = 255;
assign img[ 1798] = 255;
assign img[ 1799] = 255;
assign img[ 1800] = 255;
assign img[ 1801] = 255;
assign img[ 1802] = 255;
assign img[ 1803] = 255;
assign img[ 1804] = 255;
assign img[ 1805] = 255;
assign img[ 1806] = 255;
assign img[ 1807] = 255;
assign img[ 1808] = 255;
assign img[ 1809] = 255;
assign img[ 1810] = 255;
assign img[ 1811] = 255;
assign img[ 1812] = 255;
assign img[ 1813] = 255;
assign img[ 1814] = 255;
assign img[ 1815] = 255;
assign img[ 1816] = 255;
assign img[ 1817] = 255;
assign img[ 1818] = 255;
assign img[ 1819] = 255;
assign img[ 1820] = 255;
assign img[ 1821] = 255;
assign img[ 1822] = 255;
assign img[ 1823] = 255;
assign img[ 1824] = 255;
assign img[ 1825] = 255;
assign img[ 1826] = 255;
assign img[ 1827] = 255;
assign img[ 1828] = 255;
assign img[ 1829] = 255;
assign img[ 1830] = 255;
assign img[ 1831] = 255;
assign img[ 1832] = 255;
assign img[ 1833] = 255;
assign img[ 1834] = 255;
assign img[ 1835] = 255;
assign img[ 1836] = 255;
assign img[ 1837] = 255;
assign img[ 1838] = 255;
assign img[ 1839] = 255;
assign img[ 1840] = 255;
assign img[ 1841] = 255;
assign img[ 1842] = 255;
assign img[ 1843] = 255;
assign img[ 1844] = 255;
assign img[ 1845] = 255;
assign img[ 1846] = 255;
assign img[ 1847] = 255;
assign img[ 1848] = 255;
assign img[ 1849] = 255;
assign img[ 1850] = 255;
assign img[ 1851] = 255;
assign img[ 1852] = 255;
assign img[ 1853] = 255;
assign img[ 1854] = 255;
assign img[ 1855] = 255;
assign img[ 1856] = 255;
assign img[ 1857] = 255;
assign img[ 1858] = 255;
assign img[ 1859] = 255;
assign img[ 1860] = 255;
assign img[ 1861] = 255;
assign img[ 1862] = 255;
assign img[ 1863] = 255;
assign img[ 1864] = 255;
assign img[ 1865] = 255;
assign img[ 1866] = 255;
assign img[ 1867] = 255;
assign img[ 1868] = 255;
assign img[ 1869] = 255;
assign img[ 1870] = 255;
assign img[ 1871] = 255;
assign img[ 1872] = 255;
assign img[ 1873] = 255;
assign img[ 1874] = 255;
assign img[ 1875] = 255;
assign img[ 1876] = 255;
assign img[ 1877] = 255;
assign img[ 1878] = 255;
assign img[ 1879] = 255;
assign img[ 1880] = 255;
assign img[ 1881] = 255;
assign img[ 1882] = 255;
assign img[ 1883] = 255;
assign img[ 1884] = 255;
assign img[ 1885] = 255;
assign img[ 1886] = 255;
assign img[ 1887] = 255;
assign img[ 1888] = 255;
assign img[ 1889] = 255;
assign img[ 1890] = 255;
assign img[ 1891] = 255;
assign img[ 1892] = 255;
assign img[ 1893] = 255;
assign img[ 1894] = 255;
assign img[ 1895] = 255;
assign img[ 1896] = 255;
assign img[ 1897] = 255;
assign img[ 1898] = 255;
assign img[ 1899] = 255;
assign img[ 1900] = 255;
assign img[ 1901] = 255;
assign img[ 1902] = 255;
assign img[ 1903] = 255;
assign img[ 1904] = 255;
assign img[ 1905] = 255;
assign img[ 1906] = 255;
assign img[ 1907] = 255;
assign img[ 1908] = 255;
assign img[ 1909] = 255;
assign img[ 1910] = 255;
assign img[ 1911] = 255;
assign img[ 1912] = 255;
assign img[ 1913] = 255;
assign img[ 1914] = 255;
assign img[ 1915] = 255;
assign img[ 1916] = 255;
assign img[ 1917] = 255;
assign img[ 1918] = 255;
assign img[ 1919] = 255;
assign img[ 1920] = 255;
assign img[ 1921] = 255;
assign img[ 1922] = 255;
assign img[ 1923] = 255;
assign img[ 1924] = 255;
assign img[ 1925] = 255;
assign img[ 1926] = 255;
assign img[ 1927] = 255;
assign img[ 1928] = 255;
assign img[ 1929] = 255;
assign img[ 1930] = 255;
assign img[ 1931] = 255;
assign img[ 1932] = 255;
assign img[ 1933] = 255;
assign img[ 1934] = 255;
assign img[ 1935] = 255;
assign img[ 1936] = 255;
assign img[ 1937] = 255;
assign img[ 1938] = 255;
assign img[ 1939] = 255;
assign img[ 1940] = 255;
assign img[ 1941] = 255;
assign img[ 1942] = 255;
assign img[ 1943] = 255;
assign img[ 1944] = 255;
assign img[ 1945] = 255;
assign img[ 1946] = 255;
assign img[ 1947] = 255;
assign img[ 1948] = 255;
assign img[ 1949] = 255;
assign img[ 1950] = 255;
assign img[ 1951] = 255;
assign img[ 1952] = 255;
assign img[ 1953] = 255;
assign img[ 1954] = 255;
assign img[ 1955] = 255;
assign img[ 1956] = 255;
assign img[ 1957] = 255;
assign img[ 1958] = 255;
assign img[ 1959] = 255;
assign img[ 1960] = 255;
assign img[ 1961] = 255;
assign img[ 1962] = 255;
assign img[ 1963] = 255;
assign img[ 1964] = 255;
assign img[ 1965] = 255;
assign img[ 1966] = 255;
assign img[ 1967] = 255;
assign img[ 1968] = 255;
assign img[ 1969] = 255;
assign img[ 1970] = 255;
assign img[ 1971] = 255;
assign img[ 1972] = 255;
assign img[ 1973] = 255;
assign img[ 1974] = 255;
assign img[ 1975] = 255;
assign img[ 1976] = 255;
assign img[ 1977] = 255;
assign img[ 1978] = 255;
assign img[ 1979] = 255;
assign img[ 1980] = 255;
assign img[ 1981] = 255;
assign img[ 1982] = 255;
assign img[ 1983] = 255;
assign img[ 1984] = 255;
assign img[ 1985] = 255;
assign img[ 1986] = 255;
assign img[ 1987] = 255;
assign img[ 1988] = 255;
assign img[ 1989] = 255;
assign img[ 1990] = 255;
assign img[ 1991] = 255;
assign img[ 1992] = 255;
assign img[ 1993] = 255;
assign img[ 1994] = 255;
assign img[ 1995] = 255;
assign img[ 1996] = 255;
assign img[ 1997] = 255;
assign img[ 1998] = 255;
assign img[ 1999] = 255;
assign img[ 2000] = 255;
assign img[ 2001] = 255;
assign img[ 2002] = 255;
assign img[ 2003] = 255;
assign img[ 2004] = 255;
assign img[ 2005] = 255;
assign img[ 2006] = 255;
assign img[ 2007] = 255;
assign img[ 2008] = 255;
assign img[ 2009] = 255;
assign img[ 2010] = 255;
assign img[ 2011] = 255;
assign img[ 2012] = 255;
assign img[ 2013] = 255;
assign img[ 2014] = 255;
assign img[ 2015] = 255;
assign img[ 2016] = 255;
assign img[ 2017] = 255;
assign img[ 2018] = 255;
assign img[ 2019] = 255;
assign img[ 2020] = 255;
assign img[ 2021] = 255;
assign img[ 2022] = 255;
assign img[ 2023] = 255;
assign img[ 2024] = 255;
assign img[ 2025] = 255;
assign img[ 2026] = 255;
assign img[ 2027] = 255;
assign img[ 2028] = 255;
assign img[ 2029] = 255;
assign img[ 2030] = 255;
assign img[ 2031] = 255;
assign img[ 2032] = 255;
assign img[ 2033] = 255;
assign img[ 2034] = 255;
assign img[ 2035] = 255;
assign img[ 2036] = 255;
assign img[ 2037] = 255;
assign img[ 2038] = 255;
assign img[ 2039] = 255;
assign img[ 2040] = 255;
assign img[ 2041] = 255;
assign img[ 2042] = 255;
assign img[ 2043] = 255;
assign img[ 2044] = 255;
assign img[ 2045] = 255;
assign img[ 2046] = 255;
assign img[ 2047] = 255;
assign img[ 2048] = 221;
assign img[ 2049] = 255;
assign img[ 2050] = 255;
assign img[ 2051] = 255;
assign img[ 2052] = 255;
assign img[ 2053] = 255;
assign img[ 2054] = 255;
assign img[ 2055] = 255;
assign img[ 2056] = 255;
assign img[ 2057] = 255;
assign img[ 2058] = 255;
assign img[ 2059] = 255;
assign img[ 2060] = 255;
assign img[ 2061] = 255;
assign img[ 2062] = 255;
assign img[ 2063] = 255;
assign img[ 2064] = 255;
assign img[ 2065] = 255;
assign img[ 2066] = 255;
assign img[ 2067] = 255;
assign img[ 2068] = 255;
assign img[ 2069] = 255;
assign img[ 2070] = 255;
assign img[ 2071] = 255;
assign img[ 2072] = 255;
assign img[ 2073] = 255;
assign img[ 2074] = 255;
assign img[ 2075] = 255;
assign img[ 2076] = 255;
assign img[ 2077] = 255;
assign img[ 2078] = 255;
assign img[ 2079] = 255;
assign img[ 2080] = 255;
assign img[ 2081] = 255;
assign img[ 2082] = 255;
assign img[ 2083] = 255;
assign img[ 2084] = 255;
assign img[ 2085] = 255;
assign img[ 2086] = 255;
assign img[ 2087] = 255;
assign img[ 2088] = 255;
assign img[ 2089] = 255;
assign img[ 2090] = 255;
assign img[ 2091] = 255;
assign img[ 2092] = 255;
assign img[ 2093] = 255;
assign img[ 2094] = 255;
assign img[ 2095] = 255;
assign img[ 2096] = 255;
assign img[ 2097] = 255;
assign img[ 2098] = 255;
assign img[ 2099] = 255;
assign img[ 2100] = 255;
assign img[ 2101] = 255;
assign img[ 2102] = 255;
assign img[ 2103] = 255;
assign img[ 2104] = 255;
assign img[ 2105] = 255;
assign img[ 2106] = 255;
assign img[ 2107] = 255;
assign img[ 2108] = 255;
assign img[ 2109] = 255;
assign img[ 2110] = 255;
assign img[ 2111] = 255;
assign img[ 2112] = 255;
assign img[ 2113] = 255;
assign img[ 2114] = 255;
assign img[ 2115] = 255;
assign img[ 2116] = 255;
assign img[ 2117] = 255;
assign img[ 2118] = 255;
assign img[ 2119] = 255;
assign img[ 2120] = 255;
assign img[ 2121] = 255;
assign img[ 2122] = 255;
assign img[ 2123] = 255;
assign img[ 2124] = 255;
assign img[ 2125] = 255;
assign img[ 2126] = 255;
assign img[ 2127] = 255;
assign img[ 2128] = 255;
assign img[ 2129] = 255;
assign img[ 2130] = 255;
assign img[ 2131] = 255;
assign img[ 2132] = 255;
assign img[ 2133] = 255;
assign img[ 2134] = 255;
assign img[ 2135] = 255;
assign img[ 2136] = 255;
assign img[ 2137] = 255;
assign img[ 2138] = 255;
assign img[ 2139] = 255;
assign img[ 2140] = 255;
assign img[ 2141] = 255;
assign img[ 2142] = 255;
assign img[ 2143] = 255;
assign img[ 2144] = 255;
assign img[ 2145] = 255;
assign img[ 2146] = 255;
assign img[ 2147] = 255;
assign img[ 2148] = 255;
assign img[ 2149] = 255;
assign img[ 2150] = 255;
assign img[ 2151] = 255;
assign img[ 2152] = 255;
assign img[ 2153] = 255;
assign img[ 2154] = 255;
assign img[ 2155] = 255;
assign img[ 2156] = 255;
assign img[ 2157] = 255;
assign img[ 2158] = 255;
assign img[ 2159] = 255;
assign img[ 2160] = 255;
assign img[ 2161] = 255;
assign img[ 2162] = 255;
assign img[ 2163] = 255;
assign img[ 2164] = 255;
assign img[ 2165] = 255;
assign img[ 2166] = 255;
assign img[ 2167] = 255;
assign img[ 2168] = 255;
assign img[ 2169] = 255;
assign img[ 2170] = 255;
assign img[ 2171] = 255;
assign img[ 2172] = 255;
assign img[ 2173] = 255;
assign img[ 2174] = 255;
assign img[ 2175] = 255;
assign img[ 2176] = 255;
assign img[ 2177] = 255;
assign img[ 2178] = 255;
assign img[ 2179] = 250;
assign img[ 2180] = 254;
assign img[ 2181] = 253;
assign img[ 2182] = 248;
assign img[ 2183] = 255;
assign img[ 2184] = 249;
assign img[ 2185] = 252;
assign img[ 2186] = 247;
assign img[ 2187] = 252;
assign img[ 2188] = 254;
assign img[ 2189] = 248;
assign img[ 2190] = 255;
assign img[ 2191] = 249;
assign img[ 2192] = 248;
assign img[ 2193] = 240;
assign img[ 2194] = 254;
assign img[ 2195] = 248;
assign img[ 2196] = 254;
assign img[ 2197] = 254;
assign img[ 2198] = 248;
assign img[ 2199] = 255;
assign img[ 2200] = 255;
assign img[ 2201] = 255;
assign img[ 2202] = 254;
assign img[ 2203] = 248;
assign img[ 2204] = 248;
assign img[ 2205] = 248;
assign img[ 2206] = 254;
assign img[ 2207] = 255;
assign img[ 2208] = 255;
assign img[ 2209] = 255;
assign img[ 2210] = 248;
assign img[ 2211] = 247;
assign img[ 2212] = 248;
assign img[ 2213] = 252;
assign img[ 2214] = 254;
assign img[ 2215] = 248;
assign img[ 2216] = 248;
assign img[ 2217] = 254;
assign img[ 2218] = 248;
assign img[ 2219] = 255;
assign img[ 2220] = 248;
assign img[ 2221] = 248;
assign img[ 2222] = 248;
assign img[ 2223] = 248;
assign img[ 2224] = 255;
assign img[ 2225] = 248;
assign img[ 2226] = 248;
assign img[ 2227] = 255;
assign img[ 2228] = 255;
assign img[ 2229] = 240;
assign img[ 2230] = 248;
assign img[ 2231] = 248;
assign img[ 2232] = 252;
assign img[ 2233] = 240;
assign img[ 2234] = 245;
assign img[ 2235] = 248;
assign img[ 2236] = 252;
assign img[ 2237] = 249;
assign img[ 2238] = 249;
assign img[ 2239] = 249;
assign img[ 2240] = 252;
assign img[ 2241] = 249;
assign img[ 2242] = 252;
assign img[ 2243] = 240;
assign img[ 2244] = 246;
assign img[ 2245] = 252;
assign img[ 2246] = 251;
assign img[ 2247] = 252;
assign img[ 2248] = 251;
assign img[ 2249] = 252;
assign img[ 2250] = 240;
assign img[ 2251] = 240;
assign img[ 2252] = 240;
assign img[ 2253] = 238;
assign img[ 2254] = 252;
assign img[ 2255] = 246;
assign img[ 2256] = 254;
assign img[ 2257] = 248;
assign img[ 2258] = 240;
assign img[ 2259] = 240;
assign img[ 2260] = 254;
assign img[ 2261] = 250;
assign img[ 2262] = 240;
assign img[ 2263] = 240;
assign img[ 2264] = 254;
assign img[ 2265] = 240;
assign img[ 2266] = 240;
assign img[ 2267] = 252;
assign img[ 2268] = 252;
assign img[ 2269] = 247;
assign img[ 2270] = 255;
assign img[ 2271] = 245;
assign img[ 2272] = 245;
assign img[ 2273] = 248;
assign img[ 2274] = 245;
assign img[ 2275] = 240;
assign img[ 2276] = 239;
assign img[ 2277] = 252;
assign img[ 2278] = 253;
assign img[ 2279] = 248;
assign img[ 2280] = 252;
assign img[ 2281] = 248;
assign img[ 2282] = 253;
assign img[ 2283] = 252;
assign img[ 2284] = 248;
assign img[ 2285] = 253;
assign img[ 2286] = 239;
assign img[ 2287] = 240;
assign img[ 2288] = 252;
assign img[ 2289] = 239;
assign img[ 2290] = 240;
assign img[ 2291] = 239;
assign img[ 2292] = 252;
assign img[ 2293] = 245;
assign img[ 2294] = 240;
assign img[ 2295] = 240;
assign img[ 2296] = 240;
assign img[ 2297] = 239;
assign img[ 2298] = 252;
assign img[ 2299] = 240;
assign img[ 2300] = 240;
assign img[ 2301] = 254;
assign img[ 2302] = 252;
assign img[ 2303] = 247;
assign img[ 2304] = 239;
assign img[ 2305] = 255;
assign img[ 2306] = 255;
assign img[ 2307] = 255;
assign img[ 2308] = 255;
assign img[ 2309] = 255;
assign img[ 2310] = 255;
assign img[ 2311] = 254;
assign img[ 2312] = 255;
assign img[ 2313] = 254;
assign img[ 2314] = 254;
assign img[ 2315] = 255;
assign img[ 2316] = 255;
assign img[ 2317] = 255;
assign img[ 2318] = 255;
assign img[ 2319] = 255;
assign img[ 2320] = 255;
assign img[ 2321] = 255;
assign img[ 2322] = 255;
assign img[ 2323] = 255;
assign img[ 2324] = 255;
assign img[ 2325] = 255;
assign img[ 2326] = 255;
assign img[ 2327] = 255;
assign img[ 2328] = 255;
assign img[ 2329] = 254;
assign img[ 2330] = 255;
assign img[ 2331] = 255;
assign img[ 2332] = 255;
assign img[ 2333] = 255;
assign img[ 2334] = 255;
assign img[ 2335] = 255;
assign img[ 2336] = 255;
assign img[ 2337] = 255;
assign img[ 2338] = 255;
assign img[ 2339] = 255;
assign img[ 2340] = 255;
assign img[ 2341] = 254;
assign img[ 2342] = 255;
assign img[ 2343] = 255;
assign img[ 2344] = 255;
assign img[ 2345] = 255;
assign img[ 2346] = 253;
assign img[ 2347] = 254;
assign img[ 2348] = 248;
assign img[ 2349] = 255;
assign img[ 2350] = 255;
assign img[ 2351] = 255;
assign img[ 2352] = 255;
assign img[ 2353] = 255;
assign img[ 2354] = 255;
assign img[ 2355] = 255;
assign img[ 2356] = 255;
assign img[ 2357] = 255;
assign img[ 2358] = 255;
assign img[ 2359] = 255;
assign img[ 2360] = 255;
assign img[ 2361] = 255;
assign img[ 2362] = 255;
assign img[ 2363] = 253;
assign img[ 2364] = 253;
assign img[ 2365] = 253;
assign img[ 2366] = 255;
assign img[ 2367] = 253;
assign img[ 2368] = 253;
assign img[ 2369] = 255;
assign img[ 2370] = 253;
assign img[ 2371] = 255;
assign img[ 2372] = 255;
assign img[ 2373] = 240;
assign img[ 2374] = 255;
assign img[ 2375] = 255;
assign img[ 2376] = 245;
assign img[ 2377] = 255;
assign img[ 2378] = 255;
assign img[ 2379] = 253;
assign img[ 2380] = 255;
assign img[ 2381] = 255;
assign img[ 2382] = 255;
assign img[ 2383] = 255;
assign img[ 2384] = 252;
assign img[ 2385] = 254;
assign img[ 2386] = 253;
assign img[ 2387] = 255;
assign img[ 2388] = 255;
assign img[ 2389] = 255;
assign img[ 2390] = 255;
assign img[ 2391] = 252;
assign img[ 2392] = 251;
assign img[ 2393] = 255;
assign img[ 2394] = 255;
assign img[ 2395] = 255;
assign img[ 2396] = 252;
assign img[ 2397] = 254;
assign img[ 2398] = 252;
assign img[ 2399] = 252;
assign img[ 2400] = 240;
assign img[ 2401] = 252;
assign img[ 2402] = 255;
assign img[ 2403] = 255;
assign img[ 2404] = 252;
assign img[ 2405] = 248;
assign img[ 2406] = 255;
assign img[ 2407] = 255;
assign img[ 2408] = 252;
assign img[ 2409] = 253;
assign img[ 2410] = 255;
assign img[ 2411] = 252;
assign img[ 2412] = 248;
assign img[ 2413] = 253;
assign img[ 2414] = 249;
assign img[ 2415] = 253;
assign img[ 2416] = 248;
assign img[ 2417] = 252;
assign img[ 2418] = 249;
assign img[ 2419] = 252;
assign img[ 2420] = 240;
assign img[ 2421] = 240;
assign img[ 2422] = 254;
assign img[ 2423] = 254;
assign img[ 2424] = 252;
assign img[ 2425] = 248;
assign img[ 2426] = 249;
assign img[ 2427] = 250;
assign img[ 2428] = 253;
assign img[ 2429] = 255;
assign img[ 2430] = 255;
assign img[ 2431] = 253;
assign img[ 2432] = 255;
assign img[ 2433] = 255;
assign img[ 2434] = 255;
assign img[ 2435] = 255;
assign img[ 2436] = 255;
assign img[ 2437] = 255;
assign img[ 2438] = 255;
assign img[ 2439] = 255;
assign img[ 2440] = 255;
assign img[ 2441] = 255;
assign img[ 2442] = 255;
assign img[ 2443] = 255;
assign img[ 2444] = 255;
assign img[ 2445] = 255;
assign img[ 2446] = 255;
assign img[ 2447] = 255;
assign img[ 2448] = 255;
assign img[ 2449] = 255;
assign img[ 2450] = 255;
assign img[ 2451] = 255;
assign img[ 2452] = 248;
assign img[ 2453] = 255;
assign img[ 2454] = 255;
assign img[ 2455] = 255;
assign img[ 2456] = 255;
assign img[ 2457] = 255;
assign img[ 2458] = 255;
assign img[ 2459] = 255;
assign img[ 2460] = 255;
assign img[ 2461] = 255;
assign img[ 2462] = 255;
assign img[ 2463] = 248;
assign img[ 2464] = 255;
assign img[ 2465] = 255;
assign img[ 2466] = 255;
assign img[ 2467] = 255;
assign img[ 2468] = 255;
assign img[ 2469] = 248;
assign img[ 2470] = 255;
assign img[ 2471] = 248;
assign img[ 2472] = 248;
assign img[ 2473] = 255;
assign img[ 2474] = 255;
assign img[ 2475] = 255;
assign img[ 2476] = 248;
assign img[ 2477] = 255;
assign img[ 2478] = 255;
assign img[ 2479] = 255;
assign img[ 2480] = 255;
assign img[ 2481] = 255;
assign img[ 2482] = 255;
assign img[ 2483] = 248;
assign img[ 2484] = 254;
assign img[ 2485] = 255;
assign img[ 2486] = 255;
assign img[ 2487] = 255;
assign img[ 2488] = 255;
assign img[ 2489] = 255;
assign img[ 2490] = 255;
assign img[ 2491] = 255;
assign img[ 2492] = 255;
assign img[ 2493] = 255;
assign img[ 2494] = 255;
assign img[ 2495] = 255;
assign img[ 2496] = 255;
assign img[ 2497] = 255;
assign img[ 2498] = 250;
assign img[ 2499] = 254;
assign img[ 2500] = 255;
assign img[ 2501] = 253;
assign img[ 2502] = 255;
assign img[ 2503] = 255;
assign img[ 2504] = 255;
assign img[ 2505] = 255;
assign img[ 2506] = 250;
assign img[ 2507] = 255;
assign img[ 2508] = 255;
assign img[ 2509] = 255;
assign img[ 2510] = 254;
assign img[ 2511] = 255;
assign img[ 2512] = 255;
assign img[ 2513] = 255;
assign img[ 2514] = 255;
assign img[ 2515] = 255;
assign img[ 2516] = 255;
assign img[ 2517] = 253;
assign img[ 2518] = 252;
assign img[ 2519] = 255;
assign img[ 2520] = 252;
assign img[ 2521] = 255;
assign img[ 2522] = 255;
assign img[ 2523] = 254;
assign img[ 2524] = 240;
assign img[ 2525] = 254;
assign img[ 2526] = 255;
assign img[ 2527] = 251;
assign img[ 2528] = 254;
assign img[ 2529] = 253;
assign img[ 2530] = 250;
assign img[ 2531] = 253;
assign img[ 2532] = 255;
assign img[ 2533] = 253;
assign img[ 2534] = 251;
assign img[ 2535] = 255;
assign img[ 2536] = 252;
assign img[ 2537] = 255;
assign img[ 2538] = 255;
assign img[ 2539] = 248;
assign img[ 2540] = 255;
assign img[ 2541] = 255;
assign img[ 2542] = 255;
assign img[ 2543] = 249;
assign img[ 2544] = 255;
assign img[ 2545] = 253;
assign img[ 2546] = 255;
assign img[ 2547] = 254;
assign img[ 2548] = 253;
assign img[ 2549] = 247;
assign img[ 2550] = 250;
assign img[ 2551] = 254;
assign img[ 2552] = 254;
assign img[ 2553] = 254;
assign img[ 2554] = 248;
assign img[ 2555] = 255;
assign img[ 2556] = 253;
assign img[ 2557] = 252;
assign img[ 2558] = 252;
assign img[ 2559] = 254;
assign img[ 2560] = 248;
assign img[ 2561] = 255;
assign img[ 2562] = 255;
assign img[ 2563] = 254;
assign img[ 2564] = 255;
assign img[ 2565] = 255;
assign img[ 2566] = 255;
assign img[ 2567] = 253;
assign img[ 2568] = 253;
assign img[ 2569] = 254;
assign img[ 2570] = 255;
assign img[ 2571] = 255;
assign img[ 2572] = 255;
assign img[ 2573] = 247;
assign img[ 2574] = 255;
assign img[ 2575] = 255;
assign img[ 2576] = 248;
assign img[ 2577] = 254;
assign img[ 2578] = 248;
assign img[ 2579] = 255;
assign img[ 2580] = 248;
assign img[ 2581] = 255;
assign img[ 2582] = 255;
assign img[ 2583] = 255;
assign img[ 2584] = 254;
assign img[ 2585] = 248;
assign img[ 2586] = 255;
assign img[ 2587] = 252;
assign img[ 2588] = 255;
assign img[ 2589] = 248;
assign img[ 2590] = 255;
assign img[ 2591] = 255;
assign img[ 2592] = 254;
assign img[ 2593] = 248;
assign img[ 2594] = 255;
assign img[ 2595] = 248;
assign img[ 2596] = 255;
assign img[ 2597] = 248;
assign img[ 2598] = 254;
assign img[ 2599] = 240;
assign img[ 2600] = 254;
assign img[ 2601] = 255;
assign img[ 2602] = 255;
assign img[ 2603] = 255;
assign img[ 2604] = 248;
assign img[ 2605] = 254;
assign img[ 2606] = 255;
assign img[ 2607] = 255;
assign img[ 2608] = 248;
assign img[ 2609] = 254;
assign img[ 2610] = 248;
assign img[ 2611] = 255;
assign img[ 2612] = 255;
assign img[ 2613] = 255;
assign img[ 2614] = 254;
assign img[ 2615] = 248;
assign img[ 2616] = 255;
assign img[ 2617] = 254;
assign img[ 2618] = 255;
assign img[ 2619] = 254;
assign img[ 2620] = 254;
assign img[ 2621] = 240;
assign img[ 2622] = 253;
assign img[ 2623] = 253;
assign img[ 2624] = 240;
assign img[ 2625] = 253;
assign img[ 2626] = 253;
assign img[ 2627] = 253;
assign img[ 2628] = 254;
assign img[ 2629] = 255;
assign img[ 2630] = 252;
assign img[ 2631] = 249;
assign img[ 2632] = 247;
assign img[ 2633] = 240;
assign img[ 2634] = 253;
assign img[ 2635] = 253;
assign img[ 2636] = 249;
assign img[ 2637] = 247;
assign img[ 2638] = 255;
assign img[ 2639] = 255;
assign img[ 2640] = 253;
assign img[ 2641] = 248;
assign img[ 2642] = 255;
assign img[ 2643] = 240;
assign img[ 2644] = 255;
assign img[ 2645] = 250;
assign img[ 2646] = 251;
assign img[ 2647] = 254;
assign img[ 2648] = 255;
assign img[ 2649] = 252;
assign img[ 2650] = 255;
assign img[ 2651] = 250;
assign img[ 2652] = 255;
assign img[ 2653] = 254;
assign img[ 2654] = 254;
assign img[ 2655] = 254;
assign img[ 2656] = 253;
assign img[ 2657] = 253;
assign img[ 2658] = 255;
assign img[ 2659] = 247;
assign img[ 2660] = 253;
assign img[ 2661] = 252;
assign img[ 2662] = 255;
assign img[ 2663] = 255;
assign img[ 2664] = 249;
assign img[ 2665] = 255;
assign img[ 2666] = 240;
assign img[ 2667] = 247;
assign img[ 2668] = 253;
assign img[ 2669] = 240;
assign img[ 2670] = 253;
assign img[ 2671] = 253;
assign img[ 2672] = 255;
assign img[ 2673] = 251;
assign img[ 2674] = 252;
assign img[ 2675] = 252;
assign img[ 2676] = 240;
assign img[ 2677] = 252;
assign img[ 2678] = 251;
assign img[ 2679] = 247;
assign img[ 2680] = 252;
assign img[ 2681] = 252;
assign img[ 2682] = 253;
assign img[ 2683] = 240;
assign img[ 2684] = 254;
assign img[ 2685] = 240;
assign img[ 2686] = 255;
assign img[ 2687] = 240;
assign img[ 2688] = 253;
assign img[ 2689] = 255;
assign img[ 2690] = 252;
assign img[ 2691] = 254;
assign img[ 2692] = 253;
assign img[ 2693] = 255;
assign img[ 2694] = 255;
assign img[ 2695] = 248;
assign img[ 2696] = 248;
assign img[ 2697] = 249;
assign img[ 2698] = 248;
assign img[ 2699] = 248;
assign img[ 2700] = 255;
assign img[ 2701] = 255;
assign img[ 2702] = 255;
assign img[ 2703] = 248;
assign img[ 2704] = 248;
assign img[ 2705] = 248;
assign img[ 2706] = 248;
assign img[ 2707] = 248;
assign img[ 2708] = 248;
assign img[ 2709] = 248;
assign img[ 2710] = 248;
assign img[ 2711] = 248;
assign img[ 2712] = 248;
assign img[ 2713] = 248;
assign img[ 2714] = 248;
assign img[ 2715] = 248;
assign img[ 2716] = 248;
assign img[ 2717] = 248;
assign img[ 2718] = 247;
assign img[ 2719] = 248;
assign img[ 2720] = 248;
assign img[ 2721] = 255;
assign img[ 2722] = 248;
assign img[ 2723] = 248;
assign img[ 2724] = 248;
assign img[ 2725] = 248;
assign img[ 2726] = 247;
assign img[ 2727] = 248;
assign img[ 2728] = 248;
assign img[ 2729] = 248;
assign img[ 2730] = 255;
assign img[ 2731] = 248;
assign img[ 2732] = 255;
assign img[ 2733] = 255;
assign img[ 2734] = 240;
assign img[ 2735] = 248;
assign img[ 2736] = 255;
assign img[ 2737] = 248;
assign img[ 2738] = 248;
assign img[ 2739] = 255;
assign img[ 2740] = 247;
assign img[ 2741] = 255;
assign img[ 2742] = 248;
assign img[ 2743] = 247;
assign img[ 2744] = 248;
assign img[ 2745] = 240;
assign img[ 2746] = 248;
assign img[ 2747] = 248;
assign img[ 2748] = 255;
assign img[ 2749] = 248;
assign img[ 2750] = 248;
assign img[ 2751] = 244;
assign img[ 2752] = 250;
assign img[ 2753] = 243;
assign img[ 2754] = 252;
assign img[ 2755] = 252;
assign img[ 2756] = 251;
assign img[ 2757] = 253;
assign img[ 2758] = 252;
assign img[ 2759] = 248;
assign img[ 2760] = 253;
assign img[ 2761] = 248;
assign img[ 2762] = 251;
assign img[ 2763] = 240;
assign img[ 2764] = 248;
assign img[ 2765] = 249;
assign img[ 2766] = 249;
assign img[ 2767] = 252;
assign img[ 2768] = 240;
assign img[ 2769] = 239;
assign img[ 2770] = 248;
assign img[ 2771] = 252;
assign img[ 2772] = 249;
assign img[ 2773] = 240;
assign img[ 2774] = 248;
assign img[ 2775] = 240;
assign img[ 2776] = 248;
assign img[ 2777] = 253;
assign img[ 2778] = 245;
assign img[ 2779] = 248;
assign img[ 2780] = 248;
assign img[ 2781] = 240;
assign img[ 2782] = 248;
assign img[ 2783] = 249;
assign img[ 2784] = 249;
assign img[ 2785] = 252;
assign img[ 2786] = 249;
assign img[ 2787] = 240;
assign img[ 2788] = 240;
assign img[ 2789] = 250;
assign img[ 2790] = 244;
assign img[ 2791] = 249;
assign img[ 2792] = 240;
assign img[ 2793] = 249;
assign img[ 2794] = 249;
assign img[ 2795] = 252;
assign img[ 2796] = 247;
assign img[ 2797] = 240;
assign img[ 2798] = 249;
assign img[ 2799] = 245;
assign img[ 2800] = 249;
assign img[ 2801] = 249;
assign img[ 2802] = 248;
assign img[ 2803] = 244;
assign img[ 2804] = 253;
assign img[ 2805] = 239;
assign img[ 2806] = 240;
assign img[ 2807] = 240;
assign img[ 2808] = 252;
assign img[ 2809] = 240;
assign img[ 2810] = 248;
assign img[ 2811] = 247;
assign img[ 2812] = 240;
assign img[ 2813] = 245;
assign img[ 2814] = 239;
assign img[ 2815] = 248;
assign img[ 2816] = 240;
assign img[ 2817] = 255;
assign img[ 2818] = 254;
assign img[ 2819] = 240;
assign img[ 2820] = 248;
assign img[ 2821] = 253;
assign img[ 2822] = 253;
assign img[ 2823] = 248;
assign img[ 2824] = 248;
assign img[ 2825] = 252;
assign img[ 2826] = 252;
assign img[ 2827] = 254;
assign img[ 2828] = 240;
assign img[ 2829] = 247;
assign img[ 2830] = 252;
assign img[ 2831] = 248;
assign img[ 2832] = 240;
assign img[ 2833] = 255;
assign img[ 2834] = 248;
assign img[ 2835] = 246;
assign img[ 2836] = 240;
assign img[ 2837] = 255;
assign img[ 2838] = 254;
assign img[ 2839] = 251;
assign img[ 2840] = 250;
assign img[ 2841] = 252;
assign img[ 2842] = 252;
assign img[ 2843] = 250;
assign img[ 2844] = 252;
assign img[ 2845] = 245;
assign img[ 2846] = 248;
assign img[ 2847] = 248;
assign img[ 2848] = 248;
assign img[ 2849] = 248;
assign img[ 2850] = 240;
assign img[ 2851] = 254;
assign img[ 2852] = 249;
assign img[ 2853] = 248;
assign img[ 2854] = 240;
assign img[ 2855] = 252;
assign img[ 2856] = 241;
assign img[ 2857] = 248;
assign img[ 2858] = 248;
assign img[ 2859] = 240;
assign img[ 2860] = 250;
assign img[ 2861] = 254;
assign img[ 2862] = 243;
assign img[ 2863] = 248;
assign img[ 2864] = 246;
assign img[ 2865] = 240;
assign img[ 2866] = 247;
assign img[ 2867] = 250;
assign img[ 2868] = 250;
assign img[ 2869] = 249;
assign img[ 2870] = 240;
assign img[ 2871] = 252;
assign img[ 2872] = 240;
assign img[ 2873] = 252;
assign img[ 2874] = 244;
assign img[ 2875] = 248;
assign img[ 2876] = 250;
assign img[ 2877] = 249;
assign img[ 2878] = 244;
assign img[ 2879] = 250;
assign img[ 2880] = 253;
assign img[ 2881] = 244;
assign img[ 2882] = 247;
assign img[ 2883] = 240;
assign img[ 2884] = 244;
assign img[ 2885] = 251;
assign img[ 2886] = 247;
assign img[ 2887] = 244;
assign img[ 2888] = 243;
assign img[ 2889] = 248;
assign img[ 2890] = 250;
assign img[ 2891] = 244;
assign img[ 2892] = 240;
assign img[ 2893] = 237;
assign img[ 2894] = 246;
assign img[ 2895] = 245;
assign img[ 2896] = 249;
assign img[ 2897] = 240;
assign img[ 2898] = 240;
assign img[ 2899] = 252;
assign img[ 2900] = 245;
assign img[ 2901] = 246;
assign img[ 2902] = 242;
assign img[ 2903] = 240;
assign img[ 2904] = 246;
assign img[ 2905] = 247;
assign img[ 2906] = 240;
assign img[ 2907] = 245;
assign img[ 2908] = 240;
assign img[ 2909] = 245;
assign img[ 2910] = 240;
assign img[ 2911] = 240;
assign img[ 2912] = 237;
assign img[ 2913] = 238;
assign img[ 2914] = 246;
assign img[ 2915] = 246;
assign img[ 2916] = 245;
assign img[ 2917] = 248;
assign img[ 2918] = 240;
assign img[ 2919] = 237;
assign img[ 2920] = 245;
assign img[ 2921] = 240;
assign img[ 2922] = 240;
assign img[ 2923] = 240;
assign img[ 2924] = 240;
assign img[ 2925] = 241;
assign img[ 2926] = 238;
assign img[ 2927] = 240;
assign img[ 2928] = 239;
assign img[ 2929] = 237;
assign img[ 2930] = 247;
assign img[ 2931] = 240;
assign img[ 2932] = 248;
assign img[ 2933] = 240;
assign img[ 2934] = 246;
assign img[ 2935] = 240;
assign img[ 2936] = 248;
assign img[ 2937] = 239;
assign img[ 2938] = 238;
assign img[ 2939] = 240;
assign img[ 2940] = 240;
assign img[ 2941] = 240;
assign img[ 2942] = 247;
assign img[ 2943] = 240;
assign img[ 2944] = 240;
assign img[ 2945] = 255;
assign img[ 2946] = 255;
assign img[ 2947] = 255;
assign img[ 2948] = 255;
assign img[ 2949] = 255;
assign img[ 2950] = 255;
assign img[ 2951] = 255;
assign img[ 2952] = 255;
assign img[ 2953] = 255;
assign img[ 2954] = 255;
assign img[ 2955] = 255;
assign img[ 2956] = 255;
assign img[ 2957] = 255;
assign img[ 2958] = 255;
assign img[ 2959] = 255;
assign img[ 2960] = 255;
assign img[ 2961] = 255;
assign img[ 2962] = 255;
assign img[ 2963] = 255;
assign img[ 2964] = 255;
assign img[ 2965] = 255;
assign img[ 2966] = 255;
assign img[ 2967] = 255;
assign img[ 2968] = 255;
assign img[ 2969] = 255;
assign img[ 2970] = 255;
assign img[ 2971] = 255;
assign img[ 2972] = 255;
assign img[ 2973] = 255;
assign img[ 2974] = 255;
assign img[ 2975] = 255;
assign img[ 2976] = 255;
assign img[ 2977] = 255;
assign img[ 2978] = 255;
assign img[ 2979] = 252;
assign img[ 2980] = 255;
assign img[ 2981] = 255;
assign img[ 2982] = 255;
assign img[ 2983] = 255;
assign img[ 2984] = 255;
assign img[ 2985] = 255;
assign img[ 2986] = 255;
assign img[ 2987] = 255;
assign img[ 2988] = 255;
assign img[ 2989] = 255;
assign img[ 2990] = 255;
assign img[ 2991] = 255;
assign img[ 2992] = 255;
assign img[ 2993] = 254;
assign img[ 2994] = 255;
assign img[ 2995] = 255;
assign img[ 2996] = 255;
assign img[ 2997] = 255;
assign img[ 2998] = 255;
assign img[ 2999] = 255;
assign img[ 3000] = 255;
assign img[ 3001] = 255;
assign img[ 3002] = 255;
assign img[ 3003] = 255;
assign img[ 3004] = 255;
assign img[ 3005] = 255;
assign img[ 3006] = 255;
assign img[ 3007] = 255;
assign img[ 3008] = 255;
assign img[ 3009] = 255;
assign img[ 3010] = 255;
assign img[ 3011] = 255;
assign img[ 3012] = 253;
assign img[ 3013] = 255;
assign img[ 3014] = 255;
assign img[ 3015] = 255;
assign img[ 3016] = 255;
assign img[ 3017] = 255;
assign img[ 3018] = 255;
assign img[ 3019] = 255;
assign img[ 3020] = 255;
assign img[ 3021] = 255;
assign img[ 3022] = 255;
assign img[ 3023] = 255;
assign img[ 3024] = 253;
assign img[ 3025] = 255;
assign img[ 3026] = 255;
assign img[ 3027] = 255;
assign img[ 3028] = 255;
assign img[ 3029] = 255;
assign img[ 3030] = 255;
assign img[ 3031] = 255;
assign img[ 3032] = 255;
assign img[ 3033] = 255;
assign img[ 3034] = 255;
assign img[ 3035] = 255;
assign img[ 3036] = 255;
assign img[ 3037] = 253;
assign img[ 3038] = 255;
assign img[ 3039] = 255;
assign img[ 3040] = 255;
assign img[ 3041] = 255;
assign img[ 3042] = 253;
assign img[ 3043] = 255;
assign img[ 3044] = 255;
assign img[ 3045] = 255;
assign img[ 3046] = 255;
assign img[ 3047] = 255;
assign img[ 3048] = 255;
assign img[ 3049] = 255;
assign img[ 3050] = 255;
assign img[ 3051] = 255;
assign img[ 3052] = 255;
assign img[ 3053] = 255;
assign img[ 3054] = 255;
assign img[ 3055] = 255;
assign img[ 3056] = 255;
assign img[ 3057] = 255;
assign img[ 3058] = 255;
assign img[ 3059] = 254;
assign img[ 3060] = 255;
assign img[ 3061] = 253;
assign img[ 3062] = 253;
assign img[ 3063] = 255;
assign img[ 3064] = 255;
assign img[ 3065] = 255;
assign img[ 3066] = 255;
assign img[ 3067] = 255;
assign img[ 3068] = 255;
assign img[ 3069] = 255;
assign img[ 3070] = 255;
assign img[ 3071] = 255;
assign img[ 3072] = 255;
assign img[ 3073] = 255;
assign img[ 3074] = 255;
assign img[ 3075] = 250;
assign img[ 3076] = 254;
assign img[ 3077] = 252;
assign img[ 3078] = 254;
assign img[ 3079] = 250;
assign img[ 3080] = 254;
assign img[ 3081] = 250;
assign img[ 3082] = 255;
assign img[ 3083] = 252;
assign img[ 3084] = 248;
assign img[ 3085] = 252;
assign img[ 3086] = 255;
assign img[ 3087] = 249;
assign img[ 3088] = 249;
assign img[ 3089] = 250;
assign img[ 3090] = 248;
assign img[ 3091] = 250;
assign img[ 3092] = 249;
assign img[ 3093] = 248;
assign img[ 3094] = 249;
assign img[ 3095] = 249;
assign img[ 3096] = 249;
assign img[ 3097] = 250;
assign img[ 3098] = 254;
assign img[ 3099] = 240;
assign img[ 3100] = 245;
assign img[ 3101] = 248;
assign img[ 3102] = 240;
assign img[ 3103] = 248;
assign img[ 3104] = 245;
assign img[ 3105] = 246;
assign img[ 3106] = 246;
assign img[ 3107] = 240;
assign img[ 3108] = 252;
assign img[ 3109] = 248;
assign img[ 3110] = 245;
assign img[ 3111] = 249;
assign img[ 3112] = 246;
assign img[ 3113] = 249;
assign img[ 3114] = 249;
assign img[ 3115] = 245;
assign img[ 3116] = 249;
assign img[ 3117] = 244;
assign img[ 3118] = 248;
assign img[ 3119] = 248;
assign img[ 3120] = 251;
assign img[ 3121] = 253;
assign img[ 3122] = 252;
assign img[ 3123] = 249;
assign img[ 3124] = 246;
assign img[ 3125] = 249;
assign img[ 3126] = 249;
assign img[ 3127] = 240;
assign img[ 3128] = 255;
assign img[ 3129] = 249;
assign img[ 3130] = 248;
assign img[ 3131] = 252;
assign img[ 3132] = 255;
assign img[ 3133] = 249;
assign img[ 3134] = 240;
assign img[ 3135] = 251;
assign img[ 3136] = 251;
assign img[ 3137] = 249;
assign img[ 3138] = 246;
assign img[ 3139] = 251;
assign img[ 3140] = 246;
assign img[ 3141] = 255;
assign img[ 3142] = 252;
assign img[ 3143] = 244;
assign img[ 3144] = 250;
assign img[ 3145] = 252;
assign img[ 3146] = 249;
assign img[ 3147] = 241;
assign img[ 3148] = 245;
assign img[ 3149] = 246;
assign img[ 3150] = 240;
assign img[ 3151] = 240;
assign img[ 3152] = 248;
assign img[ 3153] = 246;
assign img[ 3154] = 252;
assign img[ 3155] = 245;
assign img[ 3156] = 240;
assign img[ 3157] = 254;
assign img[ 3158] = 240;
assign img[ 3159] = 252;
assign img[ 3160] = 247;
assign img[ 3161] = 246;
assign img[ 3162] = 252;
assign img[ 3163] = 248;
assign img[ 3164] = 242;
assign img[ 3165] = 240;
assign img[ 3166] = 248;
assign img[ 3167] = 246;
assign img[ 3168] = 255;
assign img[ 3169] = 244;
assign img[ 3170] = 239;
assign img[ 3171] = 240;
assign img[ 3172] = 248;
assign img[ 3173] = 254;
assign img[ 3174] = 246;
assign img[ 3175] = 247;
assign img[ 3176] = 246;
assign img[ 3177] = 248;
assign img[ 3178] = 253;
assign img[ 3179] = 240;
assign img[ 3180] = 245;
assign img[ 3181] = 240;
assign img[ 3182] = 248;
assign img[ 3183] = 247;
assign img[ 3184] = 248;
assign img[ 3185] = 241;
assign img[ 3186] = 245;
assign img[ 3187] = 248;
assign img[ 3188] = 240;
assign img[ 3189] = 247;
assign img[ 3190] = 248;
assign img[ 3191] = 243;
assign img[ 3192] = 245;
assign img[ 3193] = 240;
assign img[ 3194] = 240;
assign img[ 3195] = 246;
assign img[ 3196] = 242;
assign img[ 3197] = 252;
assign img[ 3198] = 240;
assign img[ 3199] = 248;
assign img[ 3200] = 240;
assign img[ 3201] = 255;
assign img[ 3202] = 255;
assign img[ 3203] = 254;
assign img[ 3204] = 255;
assign img[ 3205] = 255;
assign img[ 3206] = 254;
assign img[ 3207] = 255;
assign img[ 3208] = 252;
assign img[ 3209] = 255;
assign img[ 3210] = 249;
assign img[ 3211] = 255;
assign img[ 3212] = 252;
assign img[ 3213] = 253;
assign img[ 3214] = 249;
assign img[ 3215] = 252;
assign img[ 3216] = 244;
assign img[ 3217] = 254;
assign img[ 3218] = 253;
assign img[ 3219] = 245;
assign img[ 3220] = 254;
assign img[ 3221] = 254;
assign img[ 3222] = 252;
assign img[ 3223] = 254;
assign img[ 3224] = 252;
assign img[ 3225] = 249;
assign img[ 3226] = 254;
assign img[ 3227] = 246;
assign img[ 3228] = 250;
assign img[ 3229] = 251;
assign img[ 3230] = 252;
assign img[ 3231] = 254;
assign img[ 3232] = 247;
assign img[ 3233] = 255;
assign img[ 3234] = 248;
assign img[ 3235] = 248;
assign img[ 3236] = 249;
assign img[ 3237] = 254;
assign img[ 3238] = 248;
assign img[ 3239] = 240;
assign img[ 3240] = 252;
assign img[ 3241] = 253;
assign img[ 3242] = 252;
assign img[ 3243] = 248;
assign img[ 3244] = 252;
assign img[ 3245] = 248;
assign img[ 3246] = 254;
assign img[ 3247] = 250;
assign img[ 3248] = 255;
assign img[ 3249] = 252;
assign img[ 3250] = 249;
assign img[ 3251] = 254;
assign img[ 3252] = 247;
assign img[ 3253] = 252;
assign img[ 3254] = 240;
assign img[ 3255] = 240;
assign img[ 3256] = 253;
assign img[ 3257] = 252;
assign img[ 3258] = 254;
assign img[ 3259] = 252;
assign img[ 3260] = 240;
assign img[ 3261] = 247;
assign img[ 3262] = 252;
assign img[ 3263] = 252;
assign img[ 3264] = 240;
assign img[ 3265] = 252;
assign img[ 3266] = 253;
assign img[ 3267] = 252;
assign img[ 3268] = 247;
assign img[ 3269] = 246;
assign img[ 3270] = 239;
assign img[ 3271] = 245;
assign img[ 3272] = 247;
assign img[ 3273] = 252;
assign img[ 3274] = 253;
assign img[ 3275] = 252;
assign img[ 3276] = 245;
assign img[ 3277] = 251;
assign img[ 3278] = 247;
assign img[ 3279] = 253;
assign img[ 3280] = 253;
assign img[ 3281] = 254;
assign img[ 3282] = 245;
assign img[ 3283] = 247;
assign img[ 3284] = 253;
assign img[ 3285] = 247;
assign img[ 3286] = 254;
assign img[ 3287] = 247;
assign img[ 3288] = 246;
assign img[ 3289] = 248;
assign img[ 3290] = 255;
assign img[ 3291] = 240;
assign img[ 3292] = 240;
assign img[ 3293] = 254;
assign img[ 3294] = 255;
assign img[ 3295] = 252;
assign img[ 3296] = 248;
assign img[ 3297] = 248;
assign img[ 3298] = 246;
assign img[ 3299] = 248;
assign img[ 3300] = 253;
assign img[ 3301] = 255;
assign img[ 3302] = 255;
assign img[ 3303] = 248;
assign img[ 3304] = 254;
assign img[ 3305] = 240;
assign img[ 3306] = 248;
assign img[ 3307] = 248;
assign img[ 3308] = 254;
assign img[ 3309] = 246;
assign img[ 3310] = 248;
assign img[ 3311] = 248;
assign img[ 3312] = 248;
assign img[ 3313] = 247;
assign img[ 3314] = 248;
assign img[ 3315] = 254;
assign img[ 3316] = 248;
assign img[ 3317] = 248;
assign img[ 3318] = 248;
assign img[ 3319] = 240;
assign img[ 3320] = 247;
assign img[ 3321] = 248;
assign img[ 3322] = 248;
assign img[ 3323] = 247;
assign img[ 3324] = 248;
assign img[ 3325] = 247;
assign img[ 3326] = 240;
assign img[ 3327] = 254;
assign img[ 3328] = 247;
assign img[ 3329] = 248;
assign img[ 3330] = 240;
assign img[ 3331] = 240;
assign img[ 3332] = 235;
assign img[ 3333] = 238;
assign img[ 3334] = 240;
assign img[ 3335] = 240;
assign img[ 3336] = 240;
assign img[ 3337] = 232;
assign img[ 3338] = 233;
assign img[ 3339] = 226;
assign img[ 3340] = 236;
assign img[ 3341] = 237;
assign img[ 3342] = 232;
assign img[ 3343] = 239;
assign img[ 3344] = 236;
assign img[ 3345] = 230;
assign img[ 3346] = 237;
assign img[ 3347] = 228;
assign img[ 3348] = 237;
assign img[ 3349] = 231;
assign img[ 3350] = 229;
assign img[ 3351] = 232;
assign img[ 3352] = 236;
assign img[ 3353] = 229;
assign img[ 3354] = 237;
assign img[ 3355] = 236;
assign img[ 3356] = 232;
assign img[ 3357] = 233;
assign img[ 3358] = 233;
assign img[ 3359] = 226;
assign img[ 3360] = 236;
assign img[ 3361] = 233;
assign img[ 3362] = 237;
assign img[ 3363] = 231;
assign img[ 3364] = 229;
assign img[ 3365] = 225;
assign img[ 3366] = 230;
assign img[ 3367] = 230;
assign img[ 3368] = 236;
assign img[ 3369] = 229;
assign img[ 3370] = 233;
assign img[ 3371] = 238;
assign img[ 3372] = 237;
assign img[ 3373] = 229;
assign img[ 3374] = 231;
assign img[ 3375] = 236;
assign img[ 3376] = 236;
assign img[ 3377] = 231;
assign img[ 3378] = 233;
assign img[ 3379] = 236;
assign img[ 3380] = 226;
assign img[ 3381] = 240;
assign img[ 3382] = 226;
assign img[ 3383] = 232;
assign img[ 3384] = 230;
assign img[ 3385] = 230;
assign img[ 3386] = 229;
assign img[ 3387] = 232;
assign img[ 3388] = 225;
assign img[ 3389] = 232;
assign img[ 3390] = 226;
assign img[ 3391] = 226;
assign img[ 3392] = 221;
assign img[ 3393] = 232;
assign img[ 3394] = 226;
assign img[ 3395] = 226;
assign img[ 3396] = 233;
assign img[ 3397] = 228;
assign img[ 3398] = 226;
assign img[ 3399] = 229;
assign img[ 3400] = 226;
assign img[ 3401] = 230;
assign img[ 3402] = 229;
assign img[ 3403] = 225;
assign img[ 3404] = 232;
assign img[ 3405] = 231;
assign img[ 3406] = 233;
assign img[ 3407] = 226;
assign img[ 3408] = 226;
assign img[ 3409] = 228;
assign img[ 3410] = 236;
assign img[ 3411] = 236;
assign img[ 3412] = 231;
assign img[ 3413] = 225;
assign img[ 3414] = 230;
assign img[ 3415] = 231;
assign img[ 3416] = 232;
assign img[ 3417] = 229;
assign img[ 3418] = 232;
assign img[ 3419] = 232;
assign img[ 3420] = 230;
assign img[ 3421] = 230;
assign img[ 3422] = 230;
assign img[ 3423] = 231;
assign img[ 3424] = 229;
assign img[ 3425] = 230;
assign img[ 3426] = 232;
assign img[ 3427] = 232;
assign img[ 3428] = 232;
assign img[ 3429] = 233;
assign img[ 3430] = 232;
assign img[ 3431] = 238;
assign img[ 3432] = 230;
assign img[ 3433] = 226;
assign img[ 3434] = 236;
assign img[ 3435] = 226;
assign img[ 3436] = 230;
assign img[ 3437] = 233;
assign img[ 3438] = 230;
assign img[ 3439] = 229;
assign img[ 3440] = 227;
assign img[ 3441] = 228;
assign img[ 3442] = 232;
assign img[ 3443] = 228;
assign img[ 3444] = 232;
assign img[ 3445] = 226;
assign img[ 3446] = 232;
assign img[ 3447] = 230;
assign img[ 3448] = 229;
assign img[ 3449] = 234;
assign img[ 3450] = 231;
assign img[ 3451] = 226;
assign img[ 3452] = 218;
assign img[ 3453] = 230;
assign img[ 3454] = 225;
assign img[ 3455] = 231;
assign img[ 3456] = 229;
assign img[ 3457] = 238;
assign img[ 3458] = 235;
assign img[ 3459] = 238;
assign img[ 3460] = 230;
assign img[ 3461] = 238;
assign img[ 3462] = 232;
assign img[ 3463] = 225;
assign img[ 3464] = 228;
assign img[ 3465] = 233;
assign img[ 3466] = 233;
assign img[ 3467] = 233;
assign img[ 3468] = 225;
assign img[ 3469] = 229;
assign img[ 3470] = 228;
assign img[ 3471] = 221;
assign img[ 3472] = 223;
assign img[ 3473] = 236;
assign img[ 3474] = 231;
assign img[ 3475] = 225;
assign img[ 3476] = 231;
assign img[ 3477] = 225;
assign img[ 3478] = 219;
assign img[ 3479] = 233;
assign img[ 3480] = 218;
assign img[ 3481] = 228;
assign img[ 3482] = 226;
assign img[ 3483] = 229;
assign img[ 3484] = 225;
assign img[ 3485] = 225;
assign img[ 3486] = 233;
assign img[ 3487] = 225;
assign img[ 3488] = 220;
assign img[ 3489] = 224;
assign img[ 3490] = 229;
assign img[ 3491] = 226;
assign img[ 3492] = 226;
assign img[ 3493] = 225;
assign img[ 3494] = 227;
assign img[ 3495] = 225;
assign img[ 3496] = 232;
assign img[ 3497] = 226;
assign img[ 3498] = 226;
assign img[ 3499] = 232;
assign img[ 3500] = 225;
assign img[ 3501] = 224;
assign img[ 3502] = 227;
assign img[ 3503] = 228;
assign img[ 3504] = 221;
assign img[ 3505] = 224;
assign img[ 3506] = 224;
assign img[ 3507] = 225;
assign img[ 3508] = 229;
assign img[ 3509] = 225;
assign img[ 3510] = 230;
assign img[ 3511] = 225;
assign img[ 3512] = 224;
assign img[ 3513] = 227;
assign img[ 3514] = 226;
assign img[ 3515] = 226;
assign img[ 3516] = 226;
assign img[ 3517] = 226;
assign img[ 3518] = 228;
assign img[ 3519] = 232;
assign img[ 3520] = 226;
assign img[ 3521] = 227;
assign img[ 3522] = 224;
assign img[ 3523] = 226;
assign img[ 3524] = 225;
assign img[ 3525] = 229;
assign img[ 3526] = 228;
assign img[ 3527] = 228;
assign img[ 3528] = 230;
assign img[ 3529] = 222;
assign img[ 3530] = 224;
assign img[ 3531] = 228;
assign img[ 3532] = 221;
assign img[ 3533] = 230;
assign img[ 3534] = 222;
assign img[ 3535] = 218;
assign img[ 3536] = 224;
assign img[ 3537] = 230;
assign img[ 3538] = 227;
assign img[ 3539] = 227;
assign img[ 3540] = 230;
assign img[ 3541] = 225;
assign img[ 3542] = 227;
assign img[ 3543] = 225;
assign img[ 3544] = 225;
assign img[ 3545] = 227;
assign img[ 3546] = 222;
assign img[ 3547] = 231;
assign img[ 3548] = 227;
assign img[ 3549] = 228;
assign img[ 3550] = 222;
assign img[ 3551] = 227;
assign img[ 3552] = 226;
assign img[ 3553] = 229;
assign img[ 3554] = 232;
assign img[ 3555] = 225;
assign img[ 3556] = 231;
assign img[ 3557] = 228;
assign img[ 3558] = 226;
assign img[ 3559] = 229;
assign img[ 3560] = 226;
assign img[ 3561] = 227;
assign img[ 3562] = 220;
assign img[ 3563] = 228;
assign img[ 3564] = 227;
assign img[ 3565] = 229;
assign img[ 3566] = 226;
assign img[ 3567] = 230;
assign img[ 3568] = 231;
assign img[ 3569] = 231;
assign img[ 3570] = 227;
assign img[ 3571] = 229;
assign img[ 3572] = 218;
assign img[ 3573] = 215;
assign img[ 3574] = 224;
assign img[ 3575] = 216;
assign img[ 3576] = 229;
assign img[ 3577] = 226;
assign img[ 3578] = 224;
assign img[ 3579] = 221;
assign img[ 3580] = 221;
assign img[ 3581] = 216;
assign img[ 3582] = 216;
assign img[ 3583] = 228;
assign img[ 3584] = 230;
assign img[ 3585] = 255;
assign img[ 3586] = 248;
assign img[ 3587] = 252;
assign img[ 3588] = 255;
assign img[ 3589] = 252;
assign img[ 3590] = 255;
assign img[ 3591] = 248;
assign img[ 3592] = 240;
assign img[ 3593] = 246;
assign img[ 3594] = 248;
assign img[ 3595] = 255;
assign img[ 3596] = 250;
assign img[ 3597] = 249;
assign img[ 3598] = 242;
assign img[ 3599] = 244;
assign img[ 3600] = 244;
assign img[ 3601] = 253;
assign img[ 3602] = 253;
assign img[ 3603] = 252;
assign img[ 3604] = 249;
assign img[ 3605] = 249;
assign img[ 3606] = 252;
assign img[ 3607] = 247;
assign img[ 3608] = 240;
assign img[ 3609] = 240;
assign img[ 3610] = 248;
assign img[ 3611] = 249;
assign img[ 3612] = 245;
assign img[ 3613] = 252;
assign img[ 3614] = 246;
assign img[ 3615] = 249;
assign img[ 3616] = 241;
assign img[ 3617] = 252;
assign img[ 3618] = 248;
assign img[ 3619] = 253;
assign img[ 3620] = 245;
assign img[ 3621] = 249;
assign img[ 3622] = 252;
assign img[ 3623] = 243;
assign img[ 3624] = 241;
assign img[ 3625] = 240;
assign img[ 3626] = 245;
assign img[ 3627] = 248;
assign img[ 3628] = 255;
assign img[ 3629] = 245;
assign img[ 3630] = 252;
assign img[ 3631] = 244;
assign img[ 3632] = 250;
assign img[ 3633] = 248;
assign img[ 3634] = 246;
assign img[ 3635] = 247;
assign img[ 3636] = 241;
assign img[ 3637] = 248;
assign img[ 3638] = 252;
assign img[ 3639] = 255;
assign img[ 3640] = 248;
assign img[ 3641] = 248;
assign img[ 3642] = 252;
assign img[ 3643] = 254;
assign img[ 3644] = 247;
assign img[ 3645] = 240;
assign img[ 3646] = 252;
assign img[ 3647] = 247;
assign img[ 3648] = 248;
assign img[ 3649] = 245;
assign img[ 3650] = 248;
assign img[ 3651] = 249;
assign img[ 3652] = 248;
assign img[ 3653] = 247;
assign img[ 3654] = 246;
assign img[ 3655] = 240;
assign img[ 3656] = 248;
assign img[ 3657] = 254;
assign img[ 3658] = 248;
assign img[ 3659] = 248;
assign img[ 3660] = 248;
assign img[ 3661] = 248;
assign img[ 3662] = 249;
assign img[ 3663] = 244;
assign img[ 3664] = 240;
assign img[ 3665] = 240;
assign img[ 3666] = 252;
assign img[ 3667] = 240;
assign img[ 3668] = 240;
assign img[ 3669] = 247;
assign img[ 3670] = 254;
assign img[ 3671] = 248;
assign img[ 3672] = 240;
assign img[ 3673] = 252;
assign img[ 3674] = 248;
assign img[ 3675] = 248;
assign img[ 3676] = 240;
assign img[ 3677] = 254;
assign img[ 3678] = 240;
assign img[ 3679] = 252;
assign img[ 3680] = 248;
assign img[ 3681] = 248;
assign img[ 3682] = 240;
assign img[ 3683] = 240;
assign img[ 3684] = 248;
assign img[ 3685] = 251;
assign img[ 3686] = 247;
assign img[ 3687] = 238;
assign img[ 3688] = 240;
assign img[ 3689] = 240;
assign img[ 3690] = 247;
assign img[ 3691] = 248;
assign img[ 3692] = 252;
assign img[ 3693] = 248;
assign img[ 3694] = 247;
assign img[ 3695] = 248;
assign img[ 3696] = 239;
assign img[ 3697] = 242;
assign img[ 3698] = 247;
assign img[ 3699] = 248;
assign img[ 3700] = 240;
assign img[ 3701] = 252;
assign img[ 3702] = 244;
assign img[ 3703] = 240;
assign img[ 3704] = 240;
assign img[ 3705] = 240;
assign img[ 3706] = 239;
assign img[ 3707] = 240;
assign img[ 3708] = 247;
assign img[ 3709] = 249;
assign img[ 3710] = 240;
assign img[ 3711] = 252;
assign img[ 3712] = 240;
assign img[ 3713] = 240;
assign img[ 3714] = 240;
assign img[ 3715] = 239;
assign img[ 3716] = 235;
assign img[ 3717] = 240;
assign img[ 3718] = 239;
assign img[ 3719] = 232;
assign img[ 3720] = 238;
assign img[ 3721] = 237;
assign img[ 3722] = 234;
assign img[ 3723] = 237;
assign img[ 3724] = 236;
assign img[ 3725] = 239;
assign img[ 3726] = 234;
assign img[ 3727] = 240;
assign img[ 3728] = 238;
assign img[ 3729] = 233;
assign img[ 3730] = 242;
assign img[ 3731] = 237;
assign img[ 3732] = 229;
assign img[ 3733] = 234;
assign img[ 3734] = 236;
assign img[ 3735] = 236;
assign img[ 3736] = 237;
assign img[ 3737] = 240;
assign img[ 3738] = 238;
assign img[ 3739] = 240;
assign img[ 3740] = 233;
assign img[ 3741] = 237;
assign img[ 3742] = 235;
assign img[ 3743] = 233;
assign img[ 3744] = 237;
assign img[ 3745] = 233;
assign img[ 3746] = 233;
assign img[ 3747] = 233;
assign img[ 3748] = 233;
assign img[ 3749] = 234;
assign img[ 3750] = 237;
assign img[ 3751] = 231;
assign img[ 3752] = 235;
assign img[ 3753] = 234;
assign img[ 3754] = 238;
assign img[ 3755] = 237;
assign img[ 3756] = 233;
assign img[ 3757] = 240;
assign img[ 3758] = 237;
assign img[ 3759] = 232;
assign img[ 3760] = 239;
assign img[ 3761] = 240;
assign img[ 3762] = 237;
assign img[ 3763] = 239;
assign img[ 3764] = 239;
assign img[ 3765] = 237;
assign img[ 3766] = 237;
assign img[ 3767] = 228;
assign img[ 3768] = 229;
assign img[ 3769] = 238;
assign img[ 3770] = 235;
assign img[ 3771] = 238;
assign img[ 3772] = 235;
assign img[ 3773] = 239;
assign img[ 3774] = 229;
assign img[ 3775] = 233;
assign img[ 3776] = 233;
assign img[ 3777] = 229;
assign img[ 3778] = 229;
assign img[ 3779] = 230;
assign img[ 3780] = 234;
assign img[ 3781] = 228;
assign img[ 3782] = 232;
assign img[ 3783] = 232;
assign img[ 3784] = 232;
assign img[ 3785] = 233;
assign img[ 3786] = 230;
assign img[ 3787] = 237;
assign img[ 3788] = 230;
assign img[ 3789] = 230;
assign img[ 3790] = 228;
assign img[ 3791] = 232;
assign img[ 3792] = 232;
assign img[ 3793] = 230;
assign img[ 3794] = 231;
assign img[ 3795] = 238;
assign img[ 3796] = 232;
assign img[ 3797] = 232;
assign img[ 3798] = 239;
assign img[ 3799] = 222;
assign img[ 3800] = 230;
assign img[ 3801] = 232;
assign img[ 3802] = 232;
assign img[ 3803] = 231;
assign img[ 3804] = 230;
assign img[ 3805] = 237;
assign img[ 3806] = 239;
assign img[ 3807] = 232;
assign img[ 3808] = 231;
assign img[ 3809] = 223;
assign img[ 3810] = 227;
assign img[ 3811] = 230;
assign img[ 3812] = 230;
assign img[ 3813] = 230;
assign img[ 3814] = 238;
assign img[ 3815] = 228;
assign img[ 3816] = 229;
assign img[ 3817] = 233;
assign img[ 3818] = 229;
assign img[ 3819] = 233;
assign img[ 3820] = 225;
assign img[ 3821] = 224;
assign img[ 3822] = 232;
assign img[ 3823] = 230;
assign img[ 3824] = 227;
assign img[ 3825] = 230;
assign img[ 3826] = 228;
assign img[ 3827] = 240;
assign img[ 3828] = 229;
assign img[ 3829] = 229;
assign img[ 3830] = 230;
assign img[ 3831] = 231;
assign img[ 3832] = 231;
assign img[ 3833] = 231;
assign img[ 3834] = 227;
assign img[ 3835] = 233;
assign img[ 3836] = 232;
assign img[ 3837] = 234;
assign img[ 3838] = 228;
assign img[ 3839] = 234;
assign img[ 3840] = 232;
assign img[ 3841] = 229;
assign img[ 3842] = 225;
assign img[ 3843] = 228;
assign img[ 3844] = 226;
assign img[ 3845] = 226;
assign img[ 3846] = 226;
assign img[ 3847] = 224;
assign img[ 3848] = 225;
assign img[ 3849] = 224;
assign img[ 3850] = 225;
assign img[ 3851] = 225;
assign img[ 3852] = 215;
assign img[ 3853] = 213;
assign img[ 3854] = 216;
assign img[ 3855] = 224;
assign img[ 3856] = 213;
assign img[ 3857] = 214;
assign img[ 3858] = 224;
assign img[ 3859] = 217;
assign img[ 3860] = 214;
assign img[ 3861] = 211;
assign img[ 3862] = 213;
assign img[ 3863] = 215;
assign img[ 3864] = 221;
assign img[ 3865] = 213;
assign img[ 3866] = 219;
assign img[ 3867] = 213;
assign img[ 3868] = 209;
assign img[ 3869] = 213;
assign img[ 3870] = 217;
assign img[ 3871] = 208;
assign img[ 3872] = 217;
assign img[ 3873] = 208;
assign img[ 3874] = 208;
assign img[ 3875] = 217;
assign img[ 3876] = 208;
assign img[ 3877] = 217;
assign img[ 3878] = 215;
assign img[ 3879] = 212;
assign img[ 3880] = 214;
assign img[ 3881] = 216;
assign img[ 3882] = 213;
assign img[ 3883] = 214;
assign img[ 3884] = 213;
assign img[ 3885] = 213;
assign img[ 3886] = 208;
assign img[ 3887] = 224;
assign img[ 3888] = 220;
assign img[ 3889] = 217;
assign img[ 3890] = 217;
assign img[ 3891] = 209;
assign img[ 3892] = 217;
assign img[ 3893] = 208;
assign img[ 3894] = 213;
assign img[ 3895] = 213;
assign img[ 3896] = 213;
assign img[ 3897] = 210;
assign img[ 3898] = 225;
assign img[ 3899] = 213;
assign img[ 3900] = 220;
assign img[ 3901] = 213;
assign img[ 3902] = 206;
assign img[ 3903] = 221;
assign img[ 3904] = 213;
assign img[ 3905] = 213;
assign img[ 3906] = 217;
assign img[ 3907] = 208;
assign img[ 3908] = 223;
assign img[ 3909] = 208;
assign img[ 3910] = 213;
assign img[ 3911] = 213;
assign img[ 3912] = 215;
assign img[ 3913] = 207;
assign img[ 3914] = 213;
assign img[ 3915] = 216;
assign img[ 3916] = 225;
assign img[ 3917] = 207;
assign img[ 3918] = 208;
assign img[ 3919] = 217;
assign img[ 3920] = 217;
assign img[ 3921] = 208;
assign img[ 3922] = 208;
assign img[ 3923] = 216;
assign img[ 3924] = 208;
assign img[ 3925] = 208;
assign img[ 3926] = 208;
assign img[ 3927] = 215;
assign img[ 3928] = 208;
assign img[ 3929] = 208;
assign img[ 3930] = 208;
assign img[ 3931] = 218;
assign img[ 3932] = 208;
assign img[ 3933] = 208;
assign img[ 3934] = 208;
assign img[ 3935] = 207;
assign img[ 3936] = 208;
assign img[ 3937] = 208;
assign img[ 3938] = 207;
assign img[ 3939] = 222;
assign img[ 3940] = 214;
assign img[ 3941] = 208;
assign img[ 3942] = 205;
assign img[ 3943] = 208;
assign img[ 3944] = 208;
assign img[ 3945] = 208;
assign img[ 3946] = 214;
assign img[ 3947] = 215;
assign img[ 3948] = 214;
assign img[ 3949] = 206;
assign img[ 3950] = 214;
assign img[ 3951] = 207;
assign img[ 3952] = 213;
assign img[ 3953] = 208;
assign img[ 3954] = 207;
assign img[ 3955] = 204;
assign img[ 3956] = 207;
assign img[ 3957] = 206;
assign img[ 3958] = 208;
assign img[ 3959] = 212;
assign img[ 3960] = 208;
assign img[ 3961] = 208;
assign img[ 3962] = 208;
assign img[ 3963] = 207;
assign img[ 3964] = 207;
assign img[ 3965] = 208;
assign img[ 3966] = 215;
assign img[ 3967] = 208;
assign img[ 3968] = 208;
assign img[ 3969] = 238;
assign img[ 3970] = 232;
assign img[ 3971] = 230;
assign img[ 3972] = 225;
assign img[ 3973] = 228;
assign img[ 3974] = 227;
assign img[ 3975] = 228;
assign img[ 3976] = 226;
assign img[ 3977] = 220;
assign img[ 3978] = 230;
assign img[ 3979] = 233;
assign img[ 3980] = 226;
assign img[ 3981] = 226;
assign img[ 3982] = 229;
assign img[ 3983] = 225;
assign img[ 3984] = 225;
assign img[ 3985] = 225;
assign img[ 3986] = 223;
assign img[ 3987] = 225;
assign img[ 3988] = 229;
assign img[ 3989] = 229;
assign img[ 3990] = 220;
assign img[ 3991] = 225;
assign img[ 3992] = 225;
assign img[ 3993] = 225;
assign img[ 3994] = 225;
assign img[ 3995] = 221;
assign img[ 3996] = 221;
assign img[ 3997] = 221;
assign img[ 3998] = 216;
assign img[ 3999] = 221;
assign img[ 4000] = 221;
assign img[ 4001] = 221;
assign img[ 4002] = 217;
assign img[ 4003] = 221;
assign img[ 4004] = 217;
assign img[ 4005] = 208;
assign img[ 4006] = 217;
assign img[ 4007] = 222;
assign img[ 4008] = 225;
assign img[ 4009] = 226;
assign img[ 4010] = 225;
assign img[ 4011] = 225;
assign img[ 4012] = 228;
assign img[ 4013] = 217;
assign img[ 4014] = 213;
assign img[ 4015] = 225;
assign img[ 4016] = 217;
assign img[ 4017] = 213;
assign img[ 4018] = 228;
assign img[ 4019] = 212;
assign img[ 4020] = 225;
assign img[ 4021] = 221;
assign img[ 4022] = 220;
assign img[ 4023] = 221;
assign img[ 4024] = 212;
assign img[ 4025] = 228;
assign img[ 4026] = 225;
assign img[ 4027] = 221;
assign img[ 4028] = 219;
assign img[ 4029] = 218;
assign img[ 4030] = 225;
assign img[ 4031] = 225;
assign img[ 4032] = 225;
assign img[ 4033] = 210;
assign img[ 4034] = 225;
assign img[ 4035] = 218;
assign img[ 4036] = 219;
assign img[ 4037] = 225;
assign img[ 4038] = 221;
assign img[ 4039] = 217;
assign img[ 4040] = 218;
assign img[ 4041] = 216;
assign img[ 4042] = 225;
assign img[ 4043] = 225;
assign img[ 4044] = 226;
assign img[ 4045] = 225;
assign img[ 4046] = 225;
assign img[ 4047] = 225;
assign img[ 4048] = 225;
assign img[ 4049] = 225;
assign img[ 4050] = 217;
assign img[ 4051] = 226;
assign img[ 4052] = 226;
assign img[ 4053] = 227;
assign img[ 4054] = 225;
assign img[ 4055] = 221;
assign img[ 4056] = 227;
assign img[ 4057] = 225;
assign img[ 4058] = 230;
assign img[ 4059] = 217;
assign img[ 4060] = 215;
assign img[ 4061] = 217;
assign img[ 4062] = 222;
assign img[ 4063] = 220;
assign img[ 4064] = 217;
assign img[ 4065] = 226;
assign img[ 4066] = 225;
assign img[ 4067] = 220;
assign img[ 4068] = 217;
assign img[ 4069] = 225;
assign img[ 4070] = 220;
assign img[ 4071] = 215;
assign img[ 4072] = 217;
assign img[ 4073] = 221;
assign img[ 4074] = 217;
assign img[ 4075] = 215;
assign img[ 4076] = 219;
assign img[ 4077] = 217;
assign img[ 4078] = 217;
assign img[ 4079] = 215;
assign img[ 4080] = 217;
assign img[ 4081] = 224;
assign img[ 4082] = 225;
assign img[ 4083] = 221;
assign img[ 4084] = 217;
assign img[ 4085] = 208;
assign img[ 4086] = 225;
assign img[ 4087] = 225;
assign img[ 4088] = 219;
assign img[ 4089] = 217;
assign img[ 4090] = 216;
assign img[ 4091] = 216;
assign img[ 4092] = 225;
assign img[ 4093] = 216;
assign img[ 4094] = 212;
assign img[ 4095] = 225;
assign img[ 4096] = 192;
assign img[ 4097] = 255;
assign img[ 4098] = 252;
assign img[ 4099] = 254;
assign img[ 4100] = 255;
assign img[ 4101] = 254;
assign img[ 4102] = 255;
assign img[ 4103] = 255;
assign img[ 4104] = 252;
assign img[ 4105] = 240;
assign img[ 4106] = 255;
assign img[ 4107] = 255;
assign img[ 4108] = 255;
assign img[ 4109] = 255;
assign img[ 4110] = 252;
assign img[ 4111] = 255;
assign img[ 4112] = 255;
assign img[ 4113] = 255;
assign img[ 4114] = 255;
assign img[ 4115] = 255;
assign img[ 4116] = 255;
assign img[ 4117] = 255;
assign img[ 4118] = 255;
assign img[ 4119] = 253;
assign img[ 4120] = 255;
assign img[ 4121] = 255;
assign img[ 4122] = 255;
assign img[ 4123] = 255;
assign img[ 4124] = 246;
assign img[ 4125] = 250;
assign img[ 4126] = 240;
assign img[ 4127] = 255;
assign img[ 4128] = 248;
assign img[ 4129] = 247;
assign img[ 4130] = 250;
assign img[ 4131] = 250;
assign img[ 4132] = 247;
assign img[ 4133] = 247;
assign img[ 4134] = 252;
assign img[ 4135] = 244;
assign img[ 4136] = 246;
assign img[ 4137] = 240;
assign img[ 4138] = 247;
assign img[ 4139] = 240;
assign img[ 4140] = 253;
assign img[ 4141] = 245;
assign img[ 4142] = 240;
assign img[ 4143] = 248;
assign img[ 4144] = 255;
assign img[ 4145] = 254;
assign img[ 4146] = 239;
assign img[ 4147] = 239;
assign img[ 4148] = 248;
assign img[ 4149] = 253;
assign img[ 4150] = 240;
assign img[ 4151] = 240;
assign img[ 4152] = 255;
assign img[ 4153] = 247;
assign img[ 4154] = 248;
assign img[ 4155] = 255;
assign img[ 4156] = 252;
assign img[ 4157] = 255;
assign img[ 4158] = 255;
assign img[ 4159] = 240;
assign img[ 4160] = 236;
assign img[ 4161] = 246;
assign img[ 4162] = 254;
assign img[ 4163] = 240;
assign img[ 4164] = 240;
assign img[ 4165] = 240;
assign img[ 4166] = 248;
assign img[ 4167] = 255;
assign img[ 4168] = 240;
assign img[ 4169] = 240;
assign img[ 4170] = 240;
assign img[ 4171] = 240;
assign img[ 4172] = 240;
assign img[ 4173] = 240;
assign img[ 4174] = 240;
assign img[ 4175] = 252;
assign img[ 4176] = 239;
assign img[ 4177] = 239;
assign img[ 4178] = 240;
assign img[ 4179] = 240;
assign img[ 4180] = 247;
assign img[ 4181] = 240;
assign img[ 4182] = 248;
assign img[ 4183] = 247;
assign img[ 4184] = 240;
assign img[ 4185] = 249;
assign img[ 4186] = 247;
assign img[ 4187] = 240;
assign img[ 4188] = 238;
assign img[ 4189] = 238;
assign img[ 4190] = 238;
assign img[ 4191] = 238;
assign img[ 4192] = 239;
assign img[ 4193] = 247;
assign img[ 4194] = 239;
assign img[ 4195] = 238;
assign img[ 4196] = 239;
assign img[ 4197] = 238;
assign img[ 4198] = 240;
assign img[ 4199] = 236;
assign img[ 4200] = 239;
assign img[ 4201] = 246;
assign img[ 4202] = 239;
assign img[ 4203] = 238;
assign img[ 4204] = 244;
assign img[ 4205] = 246;
assign img[ 4206] = 238;
assign img[ 4207] = 239;
assign img[ 4208] = 238;
assign img[ 4209] = 240;
assign img[ 4210] = 239;
assign img[ 4211] = 239;
assign img[ 4212] = 236;
assign img[ 4213] = 238;
assign img[ 4214] = 236;
assign img[ 4215] = 238;
assign img[ 4216] = 239;
assign img[ 4217] = 239;
assign img[ 4218] = 239;
assign img[ 4219] = 239;
assign img[ 4220] = 238;
assign img[ 4221] = 240;
assign img[ 4222] = 239;
assign img[ 4223] = 240;
assign img[ 4224] = 236;
assign img[ 4225] = 255;
assign img[ 4226] = 254;
assign img[ 4227] = 250;
assign img[ 4228] = 255;
assign img[ 4229] = 245;
assign img[ 4230] = 248;
assign img[ 4231] = 255;
assign img[ 4232] = 253;
assign img[ 4233] = 245;
assign img[ 4234] = 248;
assign img[ 4235] = 252;
assign img[ 4236] = 254;
assign img[ 4237] = 248;
assign img[ 4238] = 255;
assign img[ 4239] = 255;
assign img[ 4240] = 255;
assign img[ 4241] = 255;
assign img[ 4242] = 255;
assign img[ 4243] = 255;
assign img[ 4244] = 255;
assign img[ 4245] = 255;
assign img[ 4246] = 255;
assign img[ 4247] = 255;
assign img[ 4248] = 255;
assign img[ 4249] = 255;
assign img[ 4250] = 255;
assign img[ 4251] = 240;
assign img[ 4252] = 247;
assign img[ 4253] = 248;
assign img[ 4254] = 255;
assign img[ 4255] = 248;
assign img[ 4256] = 255;
assign img[ 4257] = 240;
assign img[ 4258] = 248;
assign img[ 4259] = 247;
assign img[ 4260] = 240;
assign img[ 4261] = 246;
assign img[ 4262] = 252;
assign img[ 4263] = 240;
assign img[ 4264] = 248;
assign img[ 4265] = 240;
assign img[ 4266] = 246;
assign img[ 4267] = 247;
assign img[ 4268] = 248;
assign img[ 4269] = 240;
assign img[ 4270] = 246;
assign img[ 4271] = 248;
assign img[ 4272] = 248;
assign img[ 4273] = 240;
assign img[ 4274] = 240;
assign img[ 4275] = 248;
assign img[ 4276] = 254;
assign img[ 4277] = 240;
assign img[ 4278] = 248;
assign img[ 4279] = 232;
assign img[ 4280] = 252;
assign img[ 4281] = 239;
assign img[ 4282] = 236;
assign img[ 4283] = 238;
assign img[ 4284] = 237;
assign img[ 4285] = 236;
assign img[ 4286] = 248;
assign img[ 4287] = 237;
assign img[ 4288] = 239;
assign img[ 4289] = 240;
assign img[ 4290] = 236;
assign img[ 4291] = 246;
assign img[ 4292] = 238;
assign img[ 4293] = 240;
assign img[ 4294] = 245;
assign img[ 4295] = 240;
assign img[ 4296] = 241;
assign img[ 4297] = 239;
assign img[ 4298] = 240;
assign img[ 4299] = 240;
assign img[ 4300] = 240;
assign img[ 4301] = 240;
assign img[ 4302] = 239;
assign img[ 4303] = 239;
assign img[ 4304] = 252;
assign img[ 4305] = 240;
assign img[ 4306] = 239;
assign img[ 4307] = 238;
assign img[ 4308] = 240;
assign img[ 4309] = 230;
assign img[ 4310] = 240;
assign img[ 4311] = 240;
assign img[ 4312] = 240;
assign img[ 4313] = 240;
assign img[ 4314] = 240;
assign img[ 4315] = 246;
assign img[ 4316] = 239;
assign img[ 4317] = 238;
assign img[ 4318] = 244;
assign img[ 4319] = 240;
assign img[ 4320] = 239;
assign img[ 4321] = 239;
assign img[ 4322] = 241;
assign img[ 4323] = 248;
assign img[ 4324] = 236;
assign img[ 4325] = 238;
assign img[ 4326] = 239;
assign img[ 4327] = 237;
assign img[ 4328] = 239;
assign img[ 4329] = 239;
assign img[ 4330] = 240;
assign img[ 4331] = 238;
assign img[ 4332] = 240;
assign img[ 4333] = 248;
assign img[ 4334] = 238;
assign img[ 4335] = 240;
assign img[ 4336] = 240;
assign img[ 4337] = 239;
assign img[ 4338] = 240;
assign img[ 4339] = 236;
assign img[ 4340] = 239;
assign img[ 4341] = 237;
assign img[ 4342] = 239;
assign img[ 4343] = 239;
assign img[ 4344] = 239;
assign img[ 4345] = 238;
assign img[ 4346] = 236;
assign img[ 4347] = 239;
assign img[ 4348] = 239;
assign img[ 4349] = 240;
assign img[ 4350] = 239;
assign img[ 4351] = 239;
assign img[ 4352] = 239;
assign img[ 4353] = 255;
assign img[ 4354] = 255;
assign img[ 4355] = 255;
assign img[ 4356] = 255;
assign img[ 4357] = 255;
assign img[ 4358] = 255;
assign img[ 4359] = 255;
assign img[ 4360] = 255;
assign img[ 4361] = 255;
assign img[ 4362] = 255;
assign img[ 4363] = 255;
assign img[ 4364] = 255;
assign img[ 4365] = 255;
assign img[ 4366] = 255;
assign img[ 4367] = 255;
assign img[ 4368] = 255;
assign img[ 4369] = 255;
assign img[ 4370] = 255;
assign img[ 4371] = 255;
assign img[ 4372] = 255;
assign img[ 4373] = 255;
assign img[ 4374] = 255;
assign img[ 4375] = 255;
assign img[ 4376] = 255;
assign img[ 4377] = 255;
assign img[ 4378] = 255;
assign img[ 4379] = 255;
assign img[ 4380] = 255;
assign img[ 4381] = 255;
assign img[ 4382] = 255;
assign img[ 4383] = 255;
assign img[ 4384] = 255;
assign img[ 4385] = 255;
assign img[ 4386] = 255;
assign img[ 4387] = 255;
assign img[ 4388] = 254;
assign img[ 4389] = 252;
assign img[ 4390] = 255;
assign img[ 4391] = 255;
assign img[ 4392] = 255;
assign img[ 4393] = 255;
assign img[ 4394] = 253;
assign img[ 4395] = 252;
assign img[ 4396] = 248;
assign img[ 4397] = 255;
assign img[ 4398] = 254;
assign img[ 4399] = 255;
assign img[ 4400] = 255;
assign img[ 4401] = 255;
assign img[ 4402] = 248;
assign img[ 4403] = 255;
assign img[ 4404] = 248;
assign img[ 4405] = 255;
assign img[ 4406] = 254;
assign img[ 4407] = 255;
assign img[ 4408] = 248;
assign img[ 4409] = 255;
assign img[ 4410] = 255;
assign img[ 4411] = 245;
assign img[ 4412] = 240;
assign img[ 4413] = 248;
assign img[ 4414] = 247;
assign img[ 4415] = 253;
assign img[ 4416] = 253;
assign img[ 4417] = 253;
assign img[ 4418] = 255;
assign img[ 4419] = 255;
assign img[ 4420] = 253;
assign img[ 4421] = 252;
assign img[ 4422] = 249;
assign img[ 4423] = 252;
assign img[ 4424] = 245;
assign img[ 4425] = 251;
assign img[ 4426] = 253;
assign img[ 4427] = 253;
assign img[ 4428] = 255;
assign img[ 4429] = 255;
assign img[ 4430] = 255;
assign img[ 4431] = 255;
assign img[ 4432] = 240;
assign img[ 4433] = 255;
assign img[ 4434] = 240;
assign img[ 4435] = 255;
assign img[ 4436] = 255;
assign img[ 4437] = 255;
assign img[ 4438] = 255;
assign img[ 4439] = 253;
assign img[ 4440] = 240;
assign img[ 4441] = 245;
assign img[ 4442] = 255;
assign img[ 4443] = 254;
assign img[ 4444] = 244;
assign img[ 4445] = 246;
assign img[ 4446] = 252;
assign img[ 4447] = 252;
assign img[ 4448] = 252;
assign img[ 4449] = 248;
assign img[ 4450] = 253;
assign img[ 4451] = 252;
assign img[ 4452] = 239;
assign img[ 4453] = 248;
assign img[ 4454] = 240;
assign img[ 4455] = 248;
assign img[ 4456] = 248;
assign img[ 4457] = 249;
assign img[ 4458] = 248;
assign img[ 4459] = 238;
assign img[ 4460] = 239;
assign img[ 4461] = 248;
assign img[ 4462] = 248;
assign img[ 4463] = 253;
assign img[ 4464] = 252;
assign img[ 4465] = 240;
assign img[ 4466] = 253;
assign img[ 4467] = 252;
assign img[ 4468] = 240;
assign img[ 4469] = 240;
assign img[ 4470] = 240;
assign img[ 4471] = 240;
assign img[ 4472] = 239;
assign img[ 4473] = 239;
assign img[ 4474] = 241;
assign img[ 4475] = 240;
assign img[ 4476] = 239;
assign img[ 4477] = 240;
assign img[ 4478] = 240;
assign img[ 4479] = 240;
assign img[ 4480] = 240;
assign img[ 4481] = 230;
assign img[ 4482] = 227;
assign img[ 4483] = 224;
assign img[ 4484] = 221;
assign img[ 4485] = 226;
assign img[ 4486] = 225;
assign img[ 4487] = 226;
assign img[ 4488] = 226;
assign img[ 4489] = 230;
assign img[ 4490] = 226;
assign img[ 4491] = 230;
assign img[ 4492] = 231;
assign img[ 4493] = 232;
assign img[ 4494] = 240;
assign img[ 4495] = 240;
assign img[ 4496] = 239;
assign img[ 4497] = 240;
assign img[ 4498] = 248;
assign img[ 4499] = 239;
assign img[ 4500] = 239;
assign img[ 4501] = 232;
assign img[ 4502] = 239;
assign img[ 4503] = 240;
assign img[ 4504] = 240;
assign img[ 4505] = 239;
assign img[ 4506] = 240;
assign img[ 4507] = 239;
assign img[ 4508] = 232;
assign img[ 4509] = 232;
assign img[ 4510] = 232;
assign img[ 4511] = 230;
assign img[ 4512] = 226;
assign img[ 4513] = 226;
assign img[ 4514] = 226;
assign img[ 4515] = 216;
assign img[ 4516] = 230;
assign img[ 4517] = 216;
assign img[ 4518] = 215;
assign img[ 4519] = 208;
assign img[ 4520] = 215;
assign img[ 4521] = 216;
assign img[ 4522] = 224;
assign img[ 4523] = 226;
assign img[ 4524] = 216;
assign img[ 4525] = 223;
assign img[ 4526] = 215;
assign img[ 4527] = 230;
assign img[ 4528] = 208;
assign img[ 4529] = 216;
assign img[ 4530] = 215;
assign img[ 4531] = 216;
assign img[ 4532] = 214;
assign img[ 4533] = 214;
assign img[ 4534] = 214;
assign img[ 4535] = 222;
assign img[ 4536] = 208;
assign img[ 4537] = 216;
assign img[ 4538] = 223;
assign img[ 4539] = 215;
assign img[ 4540] = 218;
assign img[ 4541] = 212;
assign img[ 4542] = 210;
assign img[ 4543] = 222;
assign img[ 4544] = 207;
assign img[ 4545] = 210;
assign img[ 4546] = 213;
assign img[ 4547] = 214;
assign img[ 4548] = 215;
assign img[ 4549] = 207;
assign img[ 4550] = 220;
assign img[ 4551] = 220;
assign img[ 4552] = 216;
assign img[ 4553] = 208;
assign img[ 4554] = 215;
assign img[ 4555] = 211;
assign img[ 4556] = 214;
assign img[ 4557] = 215;
assign img[ 4558] = 209;
assign img[ 4559] = 216;
assign img[ 4560] = 208;
assign img[ 4561] = 216;
assign img[ 4562] = 212;
assign img[ 4563] = 206;
assign img[ 4564] = 209;
assign img[ 4565] = 216;
assign img[ 4566] = 210;
assign img[ 4567] = 210;
assign img[ 4568] = 210;
assign img[ 4569] = 218;
assign img[ 4570] = 216;
assign img[ 4571] = 220;
assign img[ 4572] = 207;
assign img[ 4573] = 208;
assign img[ 4574] = 214;
assign img[ 4575] = 218;
assign img[ 4576] = 216;
assign img[ 4577] = 216;
assign img[ 4578] = 210;
assign img[ 4579] = 217;
assign img[ 4580] = 212;
assign img[ 4581] = 206;
assign img[ 4582] = 216;
assign img[ 4583] = 213;
assign img[ 4584] = 210;
assign img[ 4585] = 217;
assign img[ 4586] = 220;
assign img[ 4587] = 208;
assign img[ 4588] = 208;
assign img[ 4589] = 211;
assign img[ 4590] = 211;
assign img[ 4591] = 213;
assign img[ 4592] = 216;
assign img[ 4593] = 205;
assign img[ 4594] = 206;
assign img[ 4595] = 220;
assign img[ 4596] = 204;
assign img[ 4597] = 207;
assign img[ 4598] = 205;
assign img[ 4599] = 210;
assign img[ 4600] = 198;
assign img[ 4601] = 208;
assign img[ 4602] = 210;
assign img[ 4603] = 210;
assign img[ 4604] = 207;
assign img[ 4605] = 206;
assign img[ 4606] = 204;
assign img[ 4607] = 210;
assign img[ 4608] = 208;
assign img[ 4609] = 236;
assign img[ 4610] = 228;
assign img[ 4611] = 233;
assign img[ 4612] = 226;
assign img[ 4613] = 232;
assign img[ 4614] = 224;
assign img[ 4615] = 225;
assign img[ 4616] = 225;
assign img[ 4617] = 230;
assign img[ 4618] = 228;
assign img[ 4619] = 237;
assign img[ 4620] = 232;
assign img[ 4621] = 239;
assign img[ 4622] = 238;
assign img[ 4623] = 240;
assign img[ 4624] = 240;
assign img[ 4625] = 240;
assign img[ 4626] = 240;
assign img[ 4627] = 240;
assign img[ 4628] = 240;
assign img[ 4629] = 248;
assign img[ 4630] = 246;
assign img[ 4631] = 240;
assign img[ 4632] = 238;
assign img[ 4633] = 246;
assign img[ 4634] = 239;
assign img[ 4635] = 237;
assign img[ 4636] = 240;
assign img[ 4637] = 232;
assign img[ 4638] = 238;
assign img[ 4639] = 230;
assign img[ 4640] = 230;
assign img[ 4641] = 228;
assign img[ 4642] = 228;
assign img[ 4643] = 208;
assign img[ 4644] = 225;
assign img[ 4645] = 216;
assign img[ 4646] = 214;
assign img[ 4647] = 216;
assign img[ 4648] = 215;
assign img[ 4649] = 216;
assign img[ 4650] = 230;
assign img[ 4651] = 228;
assign img[ 4652] = 216;
assign img[ 4653] = 222;
assign img[ 4654] = 220;
assign img[ 4655] = 221;
assign img[ 4656] = 216;
assign img[ 4657] = 215;
assign img[ 4658] = 208;
assign img[ 4659] = 208;
assign img[ 4660] = 222;
assign img[ 4661] = 214;
assign img[ 4662] = 224;
assign img[ 4663] = 208;
assign img[ 4664] = 216;
assign img[ 4665] = 222;
assign img[ 4666] = 222;
assign img[ 4667] = 230;
assign img[ 4668] = 216;
assign img[ 4669] = 215;
assign img[ 4670] = 216;
assign img[ 4671] = 213;
assign img[ 4672] = 208;
assign img[ 4673] = 216;
assign img[ 4674] = 212;
assign img[ 4675] = 208;
assign img[ 4676] = 217;
assign img[ 4677] = 220;
assign img[ 4678] = 222;
assign img[ 4679] = 221;
assign img[ 4680] = 220;
assign img[ 4681] = 212;
assign img[ 4682] = 216;
assign img[ 4683] = 219;
assign img[ 4684] = 216;
assign img[ 4685] = 208;
assign img[ 4686] = 210;
assign img[ 4687] = 225;
assign img[ 4688] = 220;
assign img[ 4689] = 218;
assign img[ 4690] = 217;
assign img[ 4691] = 216;
assign img[ 4692] = 218;
assign img[ 4693] = 216;
assign img[ 4694] = 207;
assign img[ 4695] = 216;
assign img[ 4696] = 220;
assign img[ 4697] = 218;
assign img[ 4698] = 218;
assign img[ 4699] = 216;
assign img[ 4700] = 224;
assign img[ 4701] = 218;
assign img[ 4702] = 218;
assign img[ 4703] = 221;
assign img[ 4704] = 217;
assign img[ 4705] = 217;
assign img[ 4706] = 220;
assign img[ 4707] = 208;
assign img[ 4708] = 217;
assign img[ 4709] = 208;
assign img[ 4710] = 221;
assign img[ 4711] = 208;
assign img[ 4712] = 221;
assign img[ 4713] = 207;
assign img[ 4714] = 208;
assign img[ 4715] = 215;
assign img[ 4716] = 208;
assign img[ 4717] = 212;
assign img[ 4718] = 220;
assign img[ 4719] = 213;
assign img[ 4720] = 215;
assign img[ 4721] = 211;
assign img[ 4722] = 220;
assign img[ 4723] = 207;
assign img[ 4724] = 216;
assign img[ 4725] = 216;
assign img[ 4726] = 208;
assign img[ 4727] = 215;
assign img[ 4728] = 213;
assign img[ 4729] = 207;
assign img[ 4730] = 221;
assign img[ 4731] = 208;
assign img[ 4732] = 208;
assign img[ 4733] = 207;
assign img[ 4734] = 206;
assign img[ 4735] = 208;
assign img[ 4736] = 208;
assign img[ 4737] = 236;
assign img[ 4738] = 227;
assign img[ 4739] = 229;
assign img[ 4740] = 225;
assign img[ 4741] = 232;
assign img[ 4742] = 236;
assign img[ 4743] = 228;
assign img[ 4744] = 224;
assign img[ 4745] = 233;
assign img[ 4746] = 230;
assign img[ 4747] = 240;
assign img[ 4748] = 247;
assign img[ 4749] = 240;
assign img[ 4750] = 247;
assign img[ 4751] = 248;
assign img[ 4752] = 248;
assign img[ 4753] = 255;
assign img[ 4754] = 248;
assign img[ 4755] = 248;
assign img[ 4756] = 248;
assign img[ 4757] = 248;
assign img[ 4758] = 255;
assign img[ 4759] = 248;
assign img[ 4760] = 255;
assign img[ 4761] = 248;
assign img[ 4762] = 240;
assign img[ 4763] = 248;
assign img[ 4764] = 240;
assign img[ 4765] = 240;
assign img[ 4766] = 232;
assign img[ 4767] = 240;
assign img[ 4768] = 240;
assign img[ 4769] = 231;
assign img[ 4770] = 231;
assign img[ 4771] = 231;
assign img[ 4772] = 226;
assign img[ 4773] = 230;
assign img[ 4774] = 226;
assign img[ 4775] = 230;
assign img[ 4776] = 230;
assign img[ 4777] = 227;
assign img[ 4778] = 231;
assign img[ 4779] = 225;
assign img[ 4780] = 227;
assign img[ 4781] = 230;
assign img[ 4782] = 230;
assign img[ 4783] = 230;
assign img[ 4784] = 225;
assign img[ 4785] = 226;
assign img[ 4786] = 216;
assign img[ 4787] = 226;
assign img[ 4788] = 228;
assign img[ 4789] = 227;
assign img[ 4790] = 216;
assign img[ 4791] = 226;
assign img[ 4792] = 227;
assign img[ 4793] = 230;
assign img[ 4794] = 229;
assign img[ 4795] = 227;
assign img[ 4796] = 226;
assign img[ 4797] = 216;
assign img[ 4798] = 222;
assign img[ 4799] = 212;
assign img[ 4800] = 224;
assign img[ 4801] = 223;
assign img[ 4802] = 216;
assign img[ 4803] = 223;
assign img[ 4804] = 221;
assign img[ 4805] = 217;
assign img[ 4806] = 222;
assign img[ 4807] = 220;
assign img[ 4808] = 214;
assign img[ 4809] = 220;
assign img[ 4810] = 225;
assign img[ 4811] = 220;
assign img[ 4812] = 222;
assign img[ 4813] = 225;
assign img[ 4814] = 220;
assign img[ 4815] = 220;
assign img[ 4816] = 208;
assign img[ 4817] = 220;
assign img[ 4818] = 216;
assign img[ 4819] = 220;
assign img[ 4820] = 216;
assign img[ 4821] = 208;
assign img[ 4822] = 216;
assign img[ 4823] = 222;
assign img[ 4824] = 217;
assign img[ 4825] = 208;
assign img[ 4826] = 224;
assign img[ 4827] = 216;
assign img[ 4828] = 220;
assign img[ 4829] = 208;
assign img[ 4830] = 220;
assign img[ 4831] = 221;
assign img[ 4832] = 220;
assign img[ 4833] = 216;
assign img[ 4834] = 217;
assign img[ 4835] = 220;
assign img[ 4836] = 216;
assign img[ 4837] = 220;
assign img[ 4838] = 220;
assign img[ 4839] = 221;
assign img[ 4840] = 221;
assign img[ 4841] = 225;
assign img[ 4842] = 221;
assign img[ 4843] = 216;
assign img[ 4844] = 215;
assign img[ 4845] = 214;
assign img[ 4846] = 213;
assign img[ 4847] = 216;
assign img[ 4848] = 221;
assign img[ 4849] = 221;
assign img[ 4850] = 208;
assign img[ 4851] = 214;
assign img[ 4852] = 221;
assign img[ 4853] = 208;
assign img[ 4854] = 214;
assign img[ 4855] = 208;
assign img[ 4856] = 220;
assign img[ 4857] = 222;
assign img[ 4858] = 208;
assign img[ 4859] = 213;
assign img[ 4860] = 214;
assign img[ 4861] = 217;
assign img[ 4862] = 221;
assign img[ 4863] = 214;
assign img[ 4864] = 214;
assign img[ 4865] = 224;
assign img[ 4866] = 230;
assign img[ 4867] = 223;
assign img[ 4868] = 226;
assign img[ 4869] = 227;
assign img[ 4870] = 224;
assign img[ 4871] = 222;
assign img[ 4872] = 222;
assign img[ 4873] = 232;
assign img[ 4874] = 220;
assign img[ 4875] = 231;
assign img[ 4876] = 236;
assign img[ 4877] = 247;
assign img[ 4878] = 239;
assign img[ 4879] = 245;
assign img[ 4880] = 240;
assign img[ 4881] = 248;
assign img[ 4882] = 252;
assign img[ 4883] = 246;
assign img[ 4884] = 240;
assign img[ 4885] = 239;
assign img[ 4886] = 235;
assign img[ 4887] = 240;
assign img[ 4888] = 236;
assign img[ 4889] = 250;
assign img[ 4890] = 240;
assign img[ 4891] = 241;
assign img[ 4892] = 240;
assign img[ 4893] = 237;
assign img[ 4894] = 236;
assign img[ 4895] = 242;
assign img[ 4896] = 239;
assign img[ 4897] = 228;
assign img[ 4898] = 226;
assign img[ 4899] = 222;
assign img[ 4900] = 217;
assign img[ 4901] = 220;
assign img[ 4902] = 216;
assign img[ 4903] = 219;
assign img[ 4904] = 217;
assign img[ 4905] = 217;
assign img[ 4906] = 225;
assign img[ 4907] = 216;
assign img[ 4908] = 225;
assign img[ 4909] = 214;
assign img[ 4910] = 217;
assign img[ 4911] = 216;
assign img[ 4912] = 214;
assign img[ 4913] = 216;
assign img[ 4914] = 220;
assign img[ 4915] = 216;
assign img[ 4916] = 212;
assign img[ 4917] = 217;
assign img[ 4918] = 208;
assign img[ 4919] = 217;
assign img[ 4920] = 220;
assign img[ 4921] = 220;
assign img[ 4922] = 215;
assign img[ 4923] = 218;
assign img[ 4924] = 216;
assign img[ 4925] = 211;
assign img[ 4926] = 217;
assign img[ 4927] = 226;
assign img[ 4928] = 214;
assign img[ 4929] = 212;
assign img[ 4930] = 219;
assign img[ 4931] = 219;
assign img[ 4932] = 216;
assign img[ 4933] = 225;
assign img[ 4934] = 217;
assign img[ 4935] = 208;
assign img[ 4936] = 213;
assign img[ 4937] = 216;
assign img[ 4938] = 216;
assign img[ 4939] = 212;
assign img[ 4940] = 222;
assign img[ 4941] = 213;
assign img[ 4942] = 224;
assign img[ 4943] = 216;
assign img[ 4944] = 209;
assign img[ 4945] = 208;
assign img[ 4946] = 216;
assign img[ 4947] = 208;
assign img[ 4948] = 213;
assign img[ 4949] = 220;
assign img[ 4950] = 213;
assign img[ 4951] = 208;
assign img[ 4952] = 214;
assign img[ 4953] = 215;
assign img[ 4954] = 213;
assign img[ 4955] = 217;
assign img[ 4956] = 208;
assign img[ 4957] = 213;
assign img[ 4958] = 205;
assign img[ 4959] = 208;
assign img[ 4960] = 221;
assign img[ 4961] = 214;
assign img[ 4962] = 213;
assign img[ 4963] = 214;
assign img[ 4964] = 214;
assign img[ 4965] = 216;
assign img[ 4966] = 207;
assign img[ 4967] = 216;
assign img[ 4968] = 213;
assign img[ 4969] = 208;
assign img[ 4970] = 208;
assign img[ 4971] = 208;
assign img[ 4972] = 213;
assign img[ 4973] = 210;
assign img[ 4974] = 208;
assign img[ 4975] = 208;
assign img[ 4976] = 214;
assign img[ 4977] = 209;
assign img[ 4978] = 207;
assign img[ 4979] = 208;
assign img[ 4980] = 212;
assign img[ 4981] = 216;
assign img[ 4982] = 212;
assign img[ 4983] = 208;
assign img[ 4984] = 206;
assign img[ 4985] = 207;
assign img[ 4986] = 206;
assign img[ 4987] = 208;
assign img[ 4988] = 208;
assign img[ 4989] = 208;
assign img[ 4990] = 207;
assign img[ 4991] = 208;
assign img[ 4992] = 218;
assign img[ 4993] = 233;
assign img[ 4994] = 241;
assign img[ 4995] = 224;
assign img[ 4996] = 229;
assign img[ 4997] = 238;
assign img[ 4998] = 225;
assign img[ 4999] = 225;
assign img[ 5000] = 232;
assign img[ 5001] = 233;
assign img[ 5002] = 233;
assign img[ 5003] = 238;
assign img[ 5004] = 237;
assign img[ 5005] = 241;
assign img[ 5006] = 249;
assign img[ 5007] = 253;
assign img[ 5008] = 253;
assign img[ 5009] = 253;
assign img[ 5010] = 249;
assign img[ 5011] = 247;
assign img[ 5012] = 253;
assign img[ 5013] = 248;
assign img[ 5014] = 249;
assign img[ 5015] = 253;
assign img[ 5016] = 245;
assign img[ 5017] = 253;
assign img[ 5018] = 249;
assign img[ 5019] = 249;
assign img[ 5020] = 248;
assign img[ 5021] = 253;
assign img[ 5022] = 246;
assign img[ 5023] = 244;
assign img[ 5024] = 232;
assign img[ 5025] = 240;
assign img[ 5026] = 237;
assign img[ 5027] = 225;
assign img[ 5028] = 228;
assign img[ 5029] = 224;
assign img[ 5030] = 229;
assign img[ 5031] = 221;
assign img[ 5032] = 220;
assign img[ 5033] = 237;
assign img[ 5034] = 221;
assign img[ 5035] = 225;
assign img[ 5036] = 225;
assign img[ 5037] = 224;
assign img[ 5038] = 223;
assign img[ 5039] = 221;
assign img[ 5040] = 213;
assign img[ 5041] = 225;
assign img[ 5042] = 221;
assign img[ 5043] = 221;
assign img[ 5044] = 228;
assign img[ 5045] = 225;
assign img[ 5046] = 216;
assign img[ 5047] = 218;
assign img[ 5048] = 225;
assign img[ 5049] = 229;
assign img[ 5050] = 228;
assign img[ 5051] = 225;
assign img[ 5052] = 217;
assign img[ 5053] = 224;
assign img[ 5054] = 225;
assign img[ 5055] = 229;
assign img[ 5056] = 225;
assign img[ 5057] = 221;
assign img[ 5058] = 228;
assign img[ 5059] = 225;
assign img[ 5060] = 225;
assign img[ 5061] = 217;
assign img[ 5062] = 229;
assign img[ 5063] = 229;
assign img[ 5064] = 225;
assign img[ 5065] = 216;
assign img[ 5066] = 221;
assign img[ 5067] = 217;
assign img[ 5068] = 225;
assign img[ 5069] = 225;
assign img[ 5070] = 225;
assign img[ 5071] = 225;
assign img[ 5072] = 217;
assign img[ 5073] = 226;
assign img[ 5074] = 224;
assign img[ 5075] = 228;
assign img[ 5076] = 217;
assign img[ 5077] = 232;
assign img[ 5078] = 221;
assign img[ 5079] = 221;
assign img[ 5080] = 223;
assign img[ 5081] = 229;
assign img[ 5082] = 220;
assign img[ 5083] = 221;
assign img[ 5084] = 220;
assign img[ 5085] = 221;
assign img[ 5086] = 221;
assign img[ 5087] = 221;
assign img[ 5088] = 221;
assign img[ 5089] = 230;
assign img[ 5090] = 217;
assign img[ 5091] = 213;
assign img[ 5092] = 216;
assign img[ 5093] = 220;
assign img[ 5094] = 220;
assign img[ 5095] = 220;
assign img[ 5096] = 220;
assign img[ 5097] = 215;
assign img[ 5098] = 221;
assign img[ 5099] = 221;
assign img[ 5100] = 220;
assign img[ 5101] = 208;
assign img[ 5102] = 221;
assign img[ 5103] = 220;
assign img[ 5104] = 220;
assign img[ 5105] = 220;
assign img[ 5106] = 208;
assign img[ 5107] = 220;
assign img[ 5108] = 208;
assign img[ 5109] = 216;
assign img[ 5110] = 220;
assign img[ 5111] = 216;
assign img[ 5112] = 229;
assign img[ 5113] = 222;
assign img[ 5114] = 220;
assign img[ 5115] = 216;
assign img[ 5116] = 220;
assign img[ 5117] = 222;
assign img[ 5118] = 215;
assign img[ 5119] = 213;
assign img[ 5120] = 208;
assign img[ 5121] = 236;
assign img[ 5122] = 231;
assign img[ 5123] = 225;
assign img[ 5124] = 231;
assign img[ 5125] = 228;
assign img[ 5126] = 228;
assign img[ 5127] = 225;
assign img[ 5128] = 229;
assign img[ 5129] = 222;
assign img[ 5130] = 232;
assign img[ 5131] = 228;
assign img[ 5132] = 234;
assign img[ 5133] = 244;
assign img[ 5134] = 248;
assign img[ 5135] = 245;
assign img[ 5136] = 237;
assign img[ 5137] = 237;
assign img[ 5138] = 248;
assign img[ 5139] = 245;
assign img[ 5140] = 241;
assign img[ 5141] = 244;
assign img[ 5142] = 246;
assign img[ 5143] = 241;
assign img[ 5144] = 245;
assign img[ 5145] = 246;
assign img[ 5146] = 246;
assign img[ 5147] = 240;
assign img[ 5148] = 237;
assign img[ 5149] = 247;
assign img[ 5150] = 238;
assign img[ 5151] = 240;
assign img[ 5152] = 243;
assign img[ 5153] = 234;
assign img[ 5154] = 242;
assign img[ 5155] = 238;
assign img[ 5156] = 228;
assign img[ 5157] = 225;
assign img[ 5158] = 221;
assign img[ 5159] = 225;
assign img[ 5160] = 213;
assign img[ 5161] = 216;
assign img[ 5162] = 222;
assign img[ 5163] = 220;
assign img[ 5164] = 221;
assign img[ 5165] = 220;
assign img[ 5166] = 218;
assign img[ 5167] = 216;
assign img[ 5168] = 219;
assign img[ 5169] = 208;
assign img[ 5170] = 222;
assign img[ 5171] = 225;
assign img[ 5172] = 219;
assign img[ 5173] = 224;
assign img[ 5174] = 217;
assign img[ 5175] = 208;
assign img[ 5176] = 223;
assign img[ 5177] = 225;
assign img[ 5178] = 222;
assign img[ 5179] = 216;
assign img[ 5180] = 225;
assign img[ 5181] = 217;
assign img[ 5182] = 216;
assign img[ 5183] = 220;
assign img[ 5184] = 224;
assign img[ 5185] = 213;
assign img[ 5186] = 210;
assign img[ 5187] = 230;
assign img[ 5188] = 225;
assign img[ 5189] = 214;
assign img[ 5190] = 223;
assign img[ 5191] = 224;
assign img[ 5192] = 210;
assign img[ 5193] = 224;
assign img[ 5194] = 217;
assign img[ 5195] = 221;
assign img[ 5196] = 213;
assign img[ 5197] = 214;
assign img[ 5198] = 215;
assign img[ 5199] = 208;
assign img[ 5200] = 222;
assign img[ 5201] = 214;
assign img[ 5202] = 216;
assign img[ 5203] = 221;
assign img[ 5204] = 208;
assign img[ 5205] = 208;
assign img[ 5206] = 215;
assign img[ 5207] = 220;
assign img[ 5208] = 208;
assign img[ 5209] = 214;
assign img[ 5210] = 220;
assign img[ 5211] = 222;
assign img[ 5212] = 213;
assign img[ 5213] = 207;
assign img[ 5214] = 215;
assign img[ 5215] = 221;
assign img[ 5216] = 215;
assign img[ 5217] = 210;
assign img[ 5218] = 220;
assign img[ 5219] = 214;
assign img[ 5220] = 216;
assign img[ 5221] = 215;
assign img[ 5222] = 213;
assign img[ 5223] = 215;
assign img[ 5224] = 212;
assign img[ 5225] = 214;
assign img[ 5226] = 213;
assign img[ 5227] = 213;
assign img[ 5228] = 216;
assign img[ 5229] = 214;
assign img[ 5230] = 216;
assign img[ 5231] = 222;
assign img[ 5232] = 215;
assign img[ 5233] = 209;
assign img[ 5234] = 213;
assign img[ 5235] = 208;
assign img[ 5236] = 209;
assign img[ 5237] = 213;
assign img[ 5238] = 212;
assign img[ 5239] = 209;
assign img[ 5240] = 205;
assign img[ 5241] = 208;
assign img[ 5242] = 213;
assign img[ 5243] = 214;
assign img[ 5244] = 214;
assign img[ 5245] = 204;
assign img[ 5246] = 215;
assign img[ 5247] = 215;
assign img[ 5248] = 208;
assign img[ 5249] = 228;
assign img[ 5250] = 226;
assign img[ 5251] = 222;
assign img[ 5252] = 230;
assign img[ 5253] = 224;
assign img[ 5254] = 224;
assign img[ 5255] = 236;
assign img[ 5256] = 228;
assign img[ 5257] = 237;
assign img[ 5258] = 225;
assign img[ 5259] = 233;
assign img[ 5260] = 238;
assign img[ 5261] = 238;
assign img[ 5262] = 244;
assign img[ 5263] = 239;
assign img[ 5264] = 242;
assign img[ 5265] = 242;
assign img[ 5266] = 239;
assign img[ 5267] = 241;
assign img[ 5268] = 238;
assign img[ 5269] = 248;
assign img[ 5270] = 244;
assign img[ 5271] = 238;
assign img[ 5272] = 240;
assign img[ 5273] = 249;
assign img[ 5274] = 239;
assign img[ 5275] = 240;
assign img[ 5276] = 240;
assign img[ 5277] = 243;
assign img[ 5278] = 239;
assign img[ 5279] = 244;
assign img[ 5280] = 239;
assign img[ 5281] = 237;
assign img[ 5282] = 236;
assign img[ 5283] = 234;
assign img[ 5284] = 233;
assign img[ 5285] = 223;
assign img[ 5286] = 220;
assign img[ 5287] = 215;
assign img[ 5288] = 220;
assign img[ 5289] = 220;
assign img[ 5290] = 216;
assign img[ 5291] = 216;
assign img[ 5292] = 220;
assign img[ 5293] = 220;
assign img[ 5294] = 223;
assign img[ 5295] = 214;
assign img[ 5296] = 208;
assign img[ 5297] = 212;
assign img[ 5298] = 217;
assign img[ 5299] = 214;
assign img[ 5300] = 207;
assign img[ 5301] = 214;
assign img[ 5302] = 215;
assign img[ 5303] = 218;
assign img[ 5304] = 217;
assign img[ 5305] = 208;
assign img[ 5306] = 212;
assign img[ 5307] = 220;
assign img[ 5308] = 222;
assign img[ 5309] = 214;
assign img[ 5310] = 225;
assign img[ 5311] = 215;
assign img[ 5312] = 220;
assign img[ 5313] = 214;
assign img[ 5314] = 216;
assign img[ 5315] = 208;
assign img[ 5316] = 213;
assign img[ 5317] = 214;
assign img[ 5318] = 214;
assign img[ 5319] = 207;
assign img[ 5320] = 224;
assign img[ 5321] = 213;
assign img[ 5322] = 221;
assign img[ 5323] = 215;
assign img[ 5324] = 209;
assign img[ 5325] = 221;
assign img[ 5326] = 211;
assign img[ 5327] = 215;
assign img[ 5328] = 208;
assign img[ 5329] = 214;
assign img[ 5330] = 215;
assign img[ 5331] = 214;
assign img[ 5332] = 213;
assign img[ 5333] = 217;
assign img[ 5334] = 224;
assign img[ 5335] = 216;
assign img[ 5336] = 208;
assign img[ 5337] = 224;
assign img[ 5338] = 214;
assign img[ 5339] = 208;
assign img[ 5340] = 208;
assign img[ 5341] = 208;
assign img[ 5342] = 215;
assign img[ 5343] = 216;
assign img[ 5344] = 215;
assign img[ 5345] = 216;
assign img[ 5346] = 214;
assign img[ 5347] = 208;
assign img[ 5348] = 225;
assign img[ 5349] = 222;
assign img[ 5350] = 220;
assign img[ 5351] = 216;
assign img[ 5352] = 222;
assign img[ 5353] = 208;
assign img[ 5354] = 215;
assign img[ 5355] = 216;
assign img[ 5356] = 208;
assign img[ 5357] = 215;
assign img[ 5358] = 222;
assign img[ 5359] = 216;
assign img[ 5360] = 216;
assign img[ 5361] = 216;
assign img[ 5362] = 224;
assign img[ 5363] = 210;
assign img[ 5364] = 208;
assign img[ 5365] = 224;
assign img[ 5366] = 214;
assign img[ 5367] = 208;
assign img[ 5368] = 214;
assign img[ 5369] = 215;
assign img[ 5370] = 216;
assign img[ 5371] = 222;
assign img[ 5372] = 215;
assign img[ 5373] = 214;
assign img[ 5374] = 208;
assign img[ 5375] = 208;
assign img[ 5376] = 215;
assign img[ 5377] = 207;
assign img[ 5378] = 200;
assign img[ 5379] = 200;
assign img[ 5380] = 195;
assign img[ 5381] = 204;
assign img[ 5382] = 204;
assign img[ 5383] = 206;
assign img[ 5384] = 196;
assign img[ 5385] = 200;
assign img[ 5386] = 197;
assign img[ 5387] = 194;
assign img[ 5388] = 208;
assign img[ 5389] = 224;
assign img[ 5390] = 207;
assign img[ 5391] = 207;
assign img[ 5392] = 208;
assign img[ 5393] = 213;
assign img[ 5394] = 224;
assign img[ 5395] = 205;
assign img[ 5396] = 205;
assign img[ 5397] = 215;
assign img[ 5398] = 215;
assign img[ 5399] = 224;
assign img[ 5400] = 208;
assign img[ 5401] = 213;
assign img[ 5402] = 220;
assign img[ 5403] = 217;
assign img[ 5404] = 205;
assign img[ 5405] = 208;
assign img[ 5406] = 213;
assign img[ 5407] = 210;
assign img[ 5408] = 217;
assign img[ 5409] = 205;
assign img[ 5410] = 207;
assign img[ 5411] = 206;
assign img[ 5412] = 208;
assign img[ 5413] = 201;
assign img[ 5414] = 196;
assign img[ 5415] = 192;
assign img[ 5416] = 192;
assign img[ 5417] = 181;
assign img[ 5418] = 193;
assign img[ 5419] = 196;
assign img[ 5420] = 192;
assign img[ 5421] = 181;
assign img[ 5422] = 192;
assign img[ 5423] = 192;
assign img[ 5424] = 192;
assign img[ 5425] = 192;
assign img[ 5426] = 192;
assign img[ 5427] = 196;
assign img[ 5428] = 193;
assign img[ 5429] = 192;
assign img[ 5430] = 193;
assign img[ 5431] = 181;
assign img[ 5432] = 192;
assign img[ 5433] = 192;
assign img[ 5434] = 193;
assign img[ 5435] = 192;
assign img[ 5436] = 181;
assign img[ 5437] = 192;
assign img[ 5438] = 178;
assign img[ 5439] = 192;
assign img[ 5440] = 192;
assign img[ 5441] = 192;
assign img[ 5442] = 192;
assign img[ 5443] = 192;
assign img[ 5444] = 193;
assign img[ 5445] = 183;
assign img[ 5446] = 192;
assign img[ 5447] = 181;
assign img[ 5448] = 192;
assign img[ 5449] = 192;
assign img[ 5450] = 192;
assign img[ 5451] = 181;
assign img[ 5452] = 192;
assign img[ 5453] = 192;
assign img[ 5454] = 181;
assign img[ 5455] = 180;
assign img[ 5456] = 182;
assign img[ 5457] = 192;
assign img[ 5458] = 187;
assign img[ 5459] = 196;
assign img[ 5460] = 192;
assign img[ 5461] = 183;
assign img[ 5462] = 181;
assign img[ 5463] = 182;
assign img[ 5464] = 192;
assign img[ 5465] = 182;
assign img[ 5466] = 192;
assign img[ 5467] = 182;
assign img[ 5468] = 178;
assign img[ 5469] = 192;
assign img[ 5470] = 192;
assign img[ 5471] = 192;
assign img[ 5472] = 192;
assign img[ 5473] = 182;
assign img[ 5474] = 192;
assign img[ 5475] = 184;
assign img[ 5476] = 193;
assign img[ 5477] = 192;
assign img[ 5478] = 192;
assign img[ 5479] = 192;
assign img[ 5480] = 192;
assign img[ 5481] = 178;
assign img[ 5482] = 192;
assign img[ 5483] = 178;
assign img[ 5484] = 182;
assign img[ 5485] = 180;
assign img[ 5486] = 192;
assign img[ 5487] = 176;
assign img[ 5488] = 181;
assign img[ 5489] = 177;
assign img[ 5490] = 192;
assign img[ 5491] = 180;
assign img[ 5492] = 193;
assign img[ 5493] = 178;
assign img[ 5494] = 192;
assign img[ 5495] = 169;
assign img[ 5496] = 177;
assign img[ 5497] = 192;
assign img[ 5498] = 180;
assign img[ 5499] = 178;
assign img[ 5500] = 177;
assign img[ 5501] = 181;
assign img[ 5502] = 179;
assign img[ 5503] = 177;
assign img[ 5504] = 181;
assign img[ 5505] = 202;
assign img[ 5506] = 207;
assign img[ 5507] = 208;
assign img[ 5508] = 200;
assign img[ 5509] = 204;
assign img[ 5510] = 207;
assign img[ 5511] = 204;
assign img[ 5512] = 204;
assign img[ 5513] = 212;
assign img[ 5514] = 209;
assign img[ 5515] = 209;
assign img[ 5516] = 225;
assign img[ 5517] = 217;
assign img[ 5518] = 225;
assign img[ 5519] = 221;
assign img[ 5520] = 221;
assign img[ 5521] = 224;
assign img[ 5522] = 221;
assign img[ 5523] = 224;
assign img[ 5524] = 221;
assign img[ 5525] = 224;
assign img[ 5526] = 213;
assign img[ 5527] = 225;
assign img[ 5528] = 218;
assign img[ 5529] = 225;
assign img[ 5530] = 226;
assign img[ 5531] = 225;
assign img[ 5532] = 221;
assign img[ 5533] = 225;
assign img[ 5534] = 217;
assign img[ 5535] = 225;
assign img[ 5536] = 228;
assign img[ 5537] = 224;
assign img[ 5538] = 221;
assign img[ 5539] = 225;
assign img[ 5540] = 214;
assign img[ 5541] = 208;
assign img[ 5542] = 210;
assign img[ 5543] = 202;
assign img[ 5544] = 205;
assign img[ 5545] = 197;
assign img[ 5546] = 194;
assign img[ 5547] = 206;
assign img[ 5548] = 197;
assign img[ 5549] = 198;
assign img[ 5550] = 195;
assign img[ 5551] = 196;
assign img[ 5552] = 200;
assign img[ 5553] = 200;
assign img[ 5554] = 196;
assign img[ 5555] = 193;
assign img[ 5556] = 193;
assign img[ 5557] = 193;
assign img[ 5558] = 204;
assign img[ 5559] = 193;
assign img[ 5560] = 192;
assign img[ 5561] = 195;
assign img[ 5562] = 194;
assign img[ 5563] = 194;
assign img[ 5564] = 193;
assign img[ 5565] = 198;
assign img[ 5566] = 204;
assign img[ 5567] = 200;
assign img[ 5568] = 199;
assign img[ 5569] = 200;
assign img[ 5570] = 196;
assign img[ 5571] = 193;
assign img[ 5572] = 192;
assign img[ 5573] = 192;
assign img[ 5574] = 196;
assign img[ 5575] = 192;
assign img[ 5576] = 196;
assign img[ 5577] = 196;
assign img[ 5578] = 192;
assign img[ 5579] = 196;
assign img[ 5580] = 192;
assign img[ 5581] = 196;
assign img[ 5582] = 194;
assign img[ 5583] = 192;
assign img[ 5584] = 195;
assign img[ 5585] = 192;
assign img[ 5586] = 192;
assign img[ 5587] = 194;
assign img[ 5588] = 198;
assign img[ 5589] = 196;
assign img[ 5590] = 192;
assign img[ 5591] = 192;
assign img[ 5592] = 192;
assign img[ 5593] = 192;
assign img[ 5594] = 196;
assign img[ 5595] = 196;
assign img[ 5596] = 192;
assign img[ 5597] = 192;
assign img[ 5598] = 198;
assign img[ 5599] = 192;
assign img[ 5600] = 193;
assign img[ 5601] = 197;
assign img[ 5602] = 196;
assign img[ 5603] = 193;
assign img[ 5604] = 192;
assign img[ 5605] = 196;
assign img[ 5606] = 192;
assign img[ 5607] = 192;
assign img[ 5608] = 194;
assign img[ 5609] = 195;
assign img[ 5610] = 193;
assign img[ 5611] = 198;
assign img[ 5612] = 193;
assign img[ 5613] = 192;
assign img[ 5614] = 192;
assign img[ 5615] = 192;
assign img[ 5616] = 203;
assign img[ 5617] = 192;
assign img[ 5618] = 193;
assign img[ 5619] = 193;
assign img[ 5620] = 192;
assign img[ 5621] = 192;
assign img[ 5622] = 192;
assign img[ 5623] = 192;
assign img[ 5624] = 192;
assign img[ 5625] = 192;
assign img[ 5626] = 192;
assign img[ 5627] = 193;
assign img[ 5628] = 192;
assign img[ 5629] = 194;
assign img[ 5630] = 198;
assign img[ 5631] = 194;
assign img[ 5632] = 192;
assign img[ 5633] = 217;
assign img[ 5634] = 215;
assign img[ 5635] = 204;
assign img[ 5636] = 215;
assign img[ 5637] = 216;
assign img[ 5638] = 216;
assign img[ 5639] = 216;
assign img[ 5640] = 208;
assign img[ 5641] = 220;
assign img[ 5642] = 214;
assign img[ 5643] = 225;
assign img[ 5644] = 220;
assign img[ 5645] = 228;
assign img[ 5646] = 226;
assign img[ 5647] = 225;
assign img[ 5648] = 225;
assign img[ 5649] = 225;
assign img[ 5650] = 228;
assign img[ 5651] = 226;
assign img[ 5652] = 237;
assign img[ 5653] = 233;
assign img[ 5654] = 222;
assign img[ 5655] = 229;
assign img[ 5656] = 228;
assign img[ 5657] = 236;
assign img[ 5658] = 230;
assign img[ 5659] = 233;
assign img[ 5660] = 229;
assign img[ 5661] = 226;
assign img[ 5662] = 229;
assign img[ 5663] = 229;
assign img[ 5664] = 225;
assign img[ 5665] = 231;
assign img[ 5666] = 232;
assign img[ 5667] = 236;
assign img[ 5668] = 229;
assign img[ 5669] = 225;
assign img[ 5670] = 224;
assign img[ 5671] = 205;
assign img[ 5672] = 212;
assign img[ 5673] = 207;
assign img[ 5674] = 205;
assign img[ 5675] = 206;
assign img[ 5676] = 208;
assign img[ 5677] = 205;
assign img[ 5678] = 205;
assign img[ 5679] = 203;
assign img[ 5680] = 210;
assign img[ 5681] = 200;
assign img[ 5682] = 205;
assign img[ 5683] = 202;
assign img[ 5684] = 194;
assign img[ 5685] = 204;
assign img[ 5686] = 205;
assign img[ 5687] = 206;
assign img[ 5688] = 205;
assign img[ 5689] = 204;
assign img[ 5690] = 206;
assign img[ 5691] = 207;
assign img[ 5692] = 207;
assign img[ 5693] = 205;
assign img[ 5694] = 206;
assign img[ 5695] = 207;
assign img[ 5696] = 201;
assign img[ 5697] = 206;
assign img[ 5698] = 206;
assign img[ 5699] = 208;
assign img[ 5700] = 204;
assign img[ 5701] = 207;
assign img[ 5702] = 197;
assign img[ 5703] = 208;
assign img[ 5704] = 200;
assign img[ 5705] = 200;
assign img[ 5706] = 211;
assign img[ 5707] = 207;
assign img[ 5708] = 208;
assign img[ 5709] = 202;
assign img[ 5710] = 208;
assign img[ 5711] = 204;
assign img[ 5712] = 206;
assign img[ 5713] = 204;
assign img[ 5714] = 207;
assign img[ 5715] = 206;
assign img[ 5716] = 208;
assign img[ 5717] = 200;
assign img[ 5718] = 208;
assign img[ 5719] = 208;
assign img[ 5720] = 206;
assign img[ 5721] = 204;
assign img[ 5722] = 200;
assign img[ 5723] = 200;
assign img[ 5724] = 206;
assign img[ 5725] = 204;
assign img[ 5726] = 208;
assign img[ 5727] = 204;
assign img[ 5728] = 199;
assign img[ 5729] = 199;
assign img[ 5730] = 204;
assign img[ 5731] = 197;
assign img[ 5732] = 200;
assign img[ 5733] = 204;
assign img[ 5734] = 207;
assign img[ 5735] = 204;
assign img[ 5736] = 206;
assign img[ 5737] = 204;
assign img[ 5738] = 197;
assign img[ 5739] = 200;
assign img[ 5740] = 206;
assign img[ 5741] = 200;
assign img[ 5742] = 207;
assign img[ 5743] = 200;
assign img[ 5744] = 200;
assign img[ 5745] = 194;
assign img[ 5746] = 207;
assign img[ 5747] = 200;
assign img[ 5748] = 200;
assign img[ 5749] = 208;
assign img[ 5750] = 200;
assign img[ 5751] = 198;
assign img[ 5752] = 196;
assign img[ 5753] = 199;
assign img[ 5754] = 205;
assign img[ 5755] = 199;
assign img[ 5756] = 200;
assign img[ 5757] = 205;
assign img[ 5758] = 207;
assign img[ 5759] = 204;
assign img[ 5760] = 206;
assign img[ 5761] = 207;
assign img[ 5762] = 204;
assign img[ 5763] = 208;
assign img[ 5764] = 204;
assign img[ 5765] = 207;
assign img[ 5766] = 204;
assign img[ 5767] = 200;
assign img[ 5768] = 202;
assign img[ 5769] = 221;
assign img[ 5770] = 216;
assign img[ 5771] = 225;
assign img[ 5772] = 226;
assign img[ 5773] = 221;
assign img[ 5774] = 217;
assign img[ 5775] = 224;
assign img[ 5776] = 224;
assign img[ 5777] = 222;
assign img[ 5778] = 228;
assign img[ 5779] = 225;
assign img[ 5780] = 216;
assign img[ 5781] = 226;
assign img[ 5782] = 230;
assign img[ 5783] = 226;
assign img[ 5784] = 225;
assign img[ 5785] = 229;
assign img[ 5786] = 220;
assign img[ 5787] = 225;
assign img[ 5788] = 217;
assign img[ 5789] = 228;
assign img[ 5790] = 221;
assign img[ 5791] = 225;
assign img[ 5792] = 225;
assign img[ 5793] = 221;
assign img[ 5794] = 225;
assign img[ 5795] = 225;
assign img[ 5796] = 218;
assign img[ 5797] = 225;
assign img[ 5798] = 225;
assign img[ 5799] = 221;
assign img[ 5800] = 206;
assign img[ 5801] = 201;
assign img[ 5802] = 198;
assign img[ 5803] = 204;
assign img[ 5804] = 198;
assign img[ 5805] = 201;
assign img[ 5806] = 201;
assign img[ 5807] = 198;
assign img[ 5808] = 201;
assign img[ 5809] = 199;
assign img[ 5810] = 197;
assign img[ 5811] = 201;
assign img[ 5812] = 199;
assign img[ 5813] = 199;
assign img[ 5814] = 201;
assign img[ 5815] = 193;
assign img[ 5816] = 195;
assign img[ 5817] = 198;
assign img[ 5818] = 195;
assign img[ 5819] = 198;
assign img[ 5820] = 201;
assign img[ 5821] = 197;
assign img[ 5822] = 197;
assign img[ 5823] = 197;
assign img[ 5824] = 193;
assign img[ 5825] = 194;
assign img[ 5826] = 194;
assign img[ 5827] = 195;
assign img[ 5828] = 194;
assign img[ 5829] = 201;
assign img[ 5830] = 200;
assign img[ 5831] = 196;
assign img[ 5832] = 194;
assign img[ 5833] = 193;
assign img[ 5834] = 196;
assign img[ 5835] = 197;
assign img[ 5836] = 193;
assign img[ 5837] = 193;
assign img[ 5838] = 194;
assign img[ 5839] = 200;
assign img[ 5840] = 194;
assign img[ 5841] = 196;
assign img[ 5842] = 200;
assign img[ 5843] = 194;
assign img[ 5844] = 196;
assign img[ 5845] = 199;
assign img[ 5846] = 199;
assign img[ 5847] = 198;
assign img[ 5848] = 192;
assign img[ 5849] = 199;
assign img[ 5850] = 198;
assign img[ 5851] = 192;
assign img[ 5852] = 194;
assign img[ 5853] = 193;
assign img[ 5854] = 196;
assign img[ 5855] = 199;
assign img[ 5856] = 193;
assign img[ 5857] = 193;
assign img[ 5858] = 192;
assign img[ 5859] = 192;
assign img[ 5860] = 192;
assign img[ 5861] = 192;
assign img[ 5862] = 198;
assign img[ 5863] = 192;
assign img[ 5864] = 192;
assign img[ 5865] = 197;
assign img[ 5866] = 195;
assign img[ 5867] = 192;
assign img[ 5868] = 192;
assign img[ 5869] = 192;
assign img[ 5870] = 198;
assign img[ 5871] = 193;
assign img[ 5872] = 193;
assign img[ 5873] = 198;
assign img[ 5874] = 192;
assign img[ 5875] = 193;
assign img[ 5876] = 192;
assign img[ 5877] = 181;
assign img[ 5878] = 194;
assign img[ 5879] = 194;
assign img[ 5880] = 194;
assign img[ 5881] = 192;
assign img[ 5882] = 195;
assign img[ 5883] = 194;
assign img[ 5884] = 194;
assign img[ 5885] = 197;
assign img[ 5886] = 192;
assign img[ 5887] = 193;
assign img[ 5888] = 199;
assign img[ 5889] = 204;
assign img[ 5890] = 203;
assign img[ 5891] = 196;
assign img[ 5892] = 207;
assign img[ 5893] = 202;
assign img[ 5894] = 202;
assign img[ 5895] = 206;
assign img[ 5896] = 200;
assign img[ 5897] = 210;
assign img[ 5898] = 217;
assign img[ 5899] = 226;
assign img[ 5900] = 215;
assign img[ 5901] = 207;
assign img[ 5902] = 215;
assign img[ 5903] = 223;
assign img[ 5904] = 217;
assign img[ 5905] = 210;
assign img[ 5906] = 220;
assign img[ 5907] = 221;
assign img[ 5908] = 212;
assign img[ 5909] = 210;
assign img[ 5910] = 221;
assign img[ 5911] = 218;
assign img[ 5912] = 225;
assign img[ 5913] = 213;
assign img[ 5914] = 214;
assign img[ 5915] = 217;
assign img[ 5916] = 217;
assign img[ 5917] = 221;
assign img[ 5918] = 217;
assign img[ 5919] = 207;
assign img[ 5920] = 216;
assign img[ 5921] = 217;
assign img[ 5922] = 217;
assign img[ 5923] = 217;
assign img[ 5924] = 222;
assign img[ 5925] = 217;
assign img[ 5926] = 209;
assign img[ 5927] = 212;
assign img[ 5928] = 202;
assign img[ 5929] = 200;
assign img[ 5930] = 193;
assign img[ 5931] = 194;
assign img[ 5932] = 193;
assign img[ 5933] = 193;
assign img[ 5934] = 180;
assign img[ 5935] = 192;
assign img[ 5936] = 196;
assign img[ 5937] = 192;
assign img[ 5938] = 192;
assign img[ 5939] = 185;
assign img[ 5940] = 185;
assign img[ 5941] = 176;
assign img[ 5942] = 192;
assign img[ 5943] = 192;
assign img[ 5944] = 188;
assign img[ 5945] = 193;
assign img[ 5946] = 193;
assign img[ 5947] = 192;
assign img[ 5948] = 192;
assign img[ 5949] = 192;
assign img[ 5950] = 193;
assign img[ 5951] = 192;
assign img[ 5952] = 181;
assign img[ 5953] = 192;
assign img[ 5954] = 193;
assign img[ 5955] = 192;
assign img[ 5956] = 192;
assign img[ 5957] = 193;
assign img[ 5958] = 192;
assign img[ 5959] = 192;
assign img[ 5960] = 195;
assign img[ 5961] = 193;
assign img[ 5962] = 181;
assign img[ 5963] = 184;
assign img[ 5964] = 193;
assign img[ 5965] = 193;
assign img[ 5966] = 192;
assign img[ 5967] = 192;
assign img[ 5968] = 192;
assign img[ 5969] = 192;
assign img[ 5970] = 195;
assign img[ 5971] = 198;
assign img[ 5972] = 193;
assign img[ 5973] = 184;
assign img[ 5974] = 184;
assign img[ 5975] = 192;
assign img[ 5976] = 192;
assign img[ 5977] = 196;
assign img[ 5978] = 188;
assign img[ 5979] = 192;
assign img[ 5980] = 192;
assign img[ 5981] = 192;
assign img[ 5982] = 192;
assign img[ 5983] = 192;
assign img[ 5984] = 192;
assign img[ 5985] = 192;
assign img[ 5986] = 192;
assign img[ 5987] = 192;
assign img[ 5988] = 192;
assign img[ 5989] = 192;
assign img[ 5990] = 180;
assign img[ 5991] = 192;
assign img[ 5992] = 175;
assign img[ 5993] = 192;
assign img[ 5994] = 183;
assign img[ 5995] = 192;
assign img[ 5996] = 192;
assign img[ 5997] = 192;
assign img[ 5998] = 192;
assign img[ 5999] = 192;
assign img[ 6000] = 192;
assign img[ 6001] = 192;
assign img[ 6002] = 192;
assign img[ 6003] = 192;
assign img[ 6004] = 175;
assign img[ 6005] = 192;
assign img[ 6006] = 176;
assign img[ 6007] = 180;
assign img[ 6008] = 192;
assign img[ 6009] = 192;
assign img[ 6010] = 176;
assign img[ 6011] = 188;
assign img[ 6012] = 192;
assign img[ 6013] = 192;
assign img[ 6014] = 192;
assign img[ 6015] = 192;
assign img[ 6016] = 192;
assign img[ 6017] = 204;
assign img[ 6018] = 196;
assign img[ 6019] = 206;
assign img[ 6020] = 193;
assign img[ 6021] = 204;
assign img[ 6022] = 200;
assign img[ 6023] = 199;
assign img[ 6024] = 194;
assign img[ 6025] = 206;
assign img[ 6026] = 213;
assign img[ 6027] = 212;
assign img[ 6028] = 213;
assign img[ 6029] = 209;
assign img[ 6030] = 213;
assign img[ 6031] = 217;
assign img[ 6032] = 210;
assign img[ 6033] = 225;
assign img[ 6034] = 208;
assign img[ 6035] = 211;
assign img[ 6036] = 205;
assign img[ 6037] = 209;
assign img[ 6038] = 219;
assign img[ 6039] = 217;
assign img[ 6040] = 217;
assign img[ 6041] = 212;
assign img[ 6042] = 225;
assign img[ 6043] = 220;
assign img[ 6044] = 216;
assign img[ 6045] = 217;
assign img[ 6046] = 216;
assign img[ 6047] = 213;
assign img[ 6048] = 217;
assign img[ 6049] = 217;
assign img[ 6050] = 217;
assign img[ 6051] = 216;
assign img[ 6052] = 210;
assign img[ 6053] = 208;
assign img[ 6054] = 217;
assign img[ 6055] = 208;
assign img[ 6056] = 202;
assign img[ 6057] = 203;
assign img[ 6058] = 202;
assign img[ 6059] = 193;
assign img[ 6060] = 192;
assign img[ 6061] = 193;
assign img[ 6062] = 192;
assign img[ 6063] = 192;
assign img[ 6064] = 193;
assign img[ 6065] = 192;
assign img[ 6066] = 184;
assign img[ 6067] = 193;
assign img[ 6068] = 192;
assign img[ 6069] = 192;
assign img[ 6070] = 193;
assign img[ 6071] = 192;
assign img[ 6072] = 185;
assign img[ 6073] = 180;
assign img[ 6074] = 192;
assign img[ 6075] = 193;
assign img[ 6076] = 192;
assign img[ 6077] = 193;
assign img[ 6078] = 183;
assign img[ 6079] = 194;
assign img[ 6080] = 181;
assign img[ 6081] = 192;
assign img[ 6082] = 179;
assign img[ 6083] = 193;
assign img[ 6084] = 192;
assign img[ 6085] = 193;
assign img[ 6086] = 192;
assign img[ 6087] = 192;
assign img[ 6088] = 193;
assign img[ 6089] = 192;
assign img[ 6090] = 193;
assign img[ 6091] = 193;
assign img[ 6092] = 184;
assign img[ 6093] = 182;
assign img[ 6094] = 193;
assign img[ 6095] = 181;
assign img[ 6096] = 192;
assign img[ 6097] = 192;
assign img[ 6098] = 192;
assign img[ 6099] = 192;
assign img[ 6100] = 178;
assign img[ 6101] = 183;
assign img[ 6102] = 193;
assign img[ 6103] = 192;
assign img[ 6104] = 183;
assign img[ 6105] = 193;
assign img[ 6106] = 192;
assign img[ 6107] = 193;
assign img[ 6108] = 193;
assign img[ 6109] = 193;
assign img[ 6110] = 192;
assign img[ 6111] = 192;
assign img[ 6112] = 193;
assign img[ 6113] = 192;
assign img[ 6114] = 193;
assign img[ 6115] = 193;
assign img[ 6116] = 178;
assign img[ 6117] = 192;
assign img[ 6118] = 180;
assign img[ 6119] = 192;
assign img[ 6120] = 192;
assign img[ 6121] = 185;
assign img[ 6122] = 192;
assign img[ 6123] = 183;
assign img[ 6124] = 193;
assign img[ 6125] = 192;
assign img[ 6126] = 192;
assign img[ 6127] = 183;
assign img[ 6128] = 179;
assign img[ 6129] = 179;
assign img[ 6130] = 193;
assign img[ 6131] = 183;
assign img[ 6132] = 185;
assign img[ 6133] = 181;
assign img[ 6134] = 192;
assign img[ 6135] = 193;
assign img[ 6136] = 192;
assign img[ 6137] = 179;
assign img[ 6138] = 180;
assign img[ 6139] = 192;
assign img[ 6140] = 185;
assign img[ 6141] = 175;
assign img[ 6142] = 194;
assign img[ 6143] = 192;
assign img[ 6144] = 137;
assign img[ 6145] = 193;
assign img[ 6146] = 188;
assign img[ 6147] = 192;
assign img[ 6148] = 196;
assign img[ 6149] = 192;
assign img[ 6150] = 192;
assign img[ 6151] = 176;
assign img[ 6152] = 192;
assign img[ 6153] = 198;
assign img[ 6154] = 199;
assign img[ 6155] = 208;
assign img[ 6156] = 208;
assign img[ 6157] = 208;
assign img[ 6158] = 204;
assign img[ 6159] = 214;
assign img[ 6160] = 207;
assign img[ 6161] = 208;
assign img[ 6162] = 208;
assign img[ 6163] = 208;
assign img[ 6164] = 216;
assign img[ 6165] = 208;
assign img[ 6166] = 208;
assign img[ 6167] = 205;
assign img[ 6168] = 207;
assign img[ 6169] = 204;
assign img[ 6170] = 206;
assign img[ 6171] = 206;
assign img[ 6172] = 206;
assign img[ 6173] = 206;
assign img[ 6174] = 208;
assign img[ 6175] = 207;
assign img[ 6176] = 205;
assign img[ 6177] = 205;
assign img[ 6178] = 203;
assign img[ 6179] = 206;
assign img[ 6180] = 200;
assign img[ 6181] = 200;
assign img[ 6182] = 212;
assign img[ 6183] = 196;
assign img[ 6184] = 194;
assign img[ 6185] = 196;
assign img[ 6186] = 195;
assign img[ 6187] = 194;
assign img[ 6188] = 192;
assign img[ 6189] = 192;
assign img[ 6190] = 176;
assign img[ 6191] = 192;
assign img[ 6192] = 192;
assign img[ 6193] = 192;
assign img[ 6194] = 175;
assign img[ 6195] = 175;
assign img[ 6196] = 192;
assign img[ 6197] = 192;
assign img[ 6198] = 176;
assign img[ 6199] = 176;
assign img[ 6200] = 192;
assign img[ 6201] = 192;
assign img[ 6202] = 192;
assign img[ 6203] = 176;
assign img[ 6204] = 192;
assign img[ 6205] = 192;
assign img[ 6206] = 192;
assign img[ 6207] = 192;
assign img[ 6208] = 176;
assign img[ 6209] = 178;
assign img[ 6210] = 192;
assign img[ 6211] = 176;
assign img[ 6212] = 174;
assign img[ 6213] = 176;
assign img[ 6214] = 172;
assign img[ 6215] = 192;
assign img[ 6216] = 176;
assign img[ 6217] = 192;
assign img[ 6218] = 176;
assign img[ 6219] = 192;
assign img[ 6220] = 175;
assign img[ 6221] = 175;
assign img[ 6222] = 175;
assign img[ 6223] = 192;
assign img[ 6224] = 174;
assign img[ 6225] = 166;
assign img[ 6226] = 192;
assign img[ 6227] = 192;
assign img[ 6228] = 175;
assign img[ 6229] = 192;
assign img[ 6230] = 192;
assign img[ 6231] = 192;
assign img[ 6232] = 192;
assign img[ 6233] = 192;
assign img[ 6234] = 192;
assign img[ 6235] = 174;
assign img[ 6236] = 174;
assign img[ 6237] = 166;
assign img[ 6238] = 172;
assign img[ 6239] = 172;
assign img[ 6240] = 173;
assign img[ 6241] = 166;
assign img[ 6242] = 174;
assign img[ 6243] = 172;
assign img[ 6244] = 167;
assign img[ 6245] = 170;
assign img[ 6246] = 172;
assign img[ 6247] = 173;
assign img[ 6248] = 174;
assign img[ 6249] = 192;
assign img[ 6250] = 174;
assign img[ 6251] = 174;
assign img[ 6252] = 164;
assign img[ 6253] = 166;
assign img[ 6254] = 172;
assign img[ 6255] = 174;
assign img[ 6256] = 174;
assign img[ 6257] = 175;
assign img[ 6258] = 166;
assign img[ 6259] = 172;
assign img[ 6260] = 166;
assign img[ 6261] = 164;
assign img[ 6262] = 164;
assign img[ 6263] = 164;
assign img[ 6264] = 172;
assign img[ 6265] = 174;
assign img[ 6266] = 174;
assign img[ 6267] = 175;
assign img[ 6268] = 172;
assign img[ 6269] = 167;
assign img[ 6270] = 167;
assign img[ 6271] = 174;
assign img[ 6272] = 172;
assign img[ 6273] = 194;
assign img[ 6274] = 194;
assign img[ 6275] = 192;
assign img[ 6276] = 192;
assign img[ 6277] = 193;
assign img[ 6278] = 194;
assign img[ 6279] = 192;
assign img[ 6280] = 192;
assign img[ 6281] = 196;
assign img[ 6282] = 199;
assign img[ 6283] = 208;
assign img[ 6284] = 214;
assign img[ 6285] = 208;
assign img[ 6286] = 214;
assign img[ 6287] = 201;
assign img[ 6288] = 206;
assign img[ 6289] = 208;
assign img[ 6290] = 207;
assign img[ 6291] = 208;
assign img[ 6292] = 208;
assign img[ 6293] = 206;
assign img[ 6294] = 208;
assign img[ 6295] = 207;
assign img[ 6296] = 208;
assign img[ 6297] = 208;
assign img[ 6298] = 206;
assign img[ 6299] = 207;
assign img[ 6300] = 199;
assign img[ 6301] = 208;
assign img[ 6302] = 207;
assign img[ 6303] = 208;
assign img[ 6304] = 207;
assign img[ 6305] = 206;
assign img[ 6306] = 207;
assign img[ 6307] = 207;
assign img[ 6308] = 204;
assign img[ 6309] = 202;
assign img[ 6310] = 206;
assign img[ 6311] = 208;
assign img[ 6312] = 200;
assign img[ 6313] = 207;
assign img[ 6314] = 199;
assign img[ 6315] = 199;
assign img[ 6316] = 198;
assign img[ 6317] = 194;
assign img[ 6318] = 192;
assign img[ 6319] = 192;
assign img[ 6320] = 194;
assign img[ 6321] = 176;
assign img[ 6322] = 192;
assign img[ 6323] = 192;
assign img[ 6324] = 182;
assign img[ 6325] = 192;
assign img[ 6326] = 194;
assign img[ 6327] = 192;
assign img[ 6328] = 192;
assign img[ 6329] = 175;
assign img[ 6330] = 172;
assign img[ 6331] = 176;
assign img[ 6332] = 174;
assign img[ 6333] = 179;
assign img[ 6334] = 173;
assign img[ 6335] = 177;
assign img[ 6336] = 174;
assign img[ 6337] = 176;
assign img[ 6338] = 172;
assign img[ 6339] = 174;
assign img[ 6340] = 172;
assign img[ 6341] = 175;
assign img[ 6342] = 181;
assign img[ 6343] = 172;
assign img[ 6344] = 173;
assign img[ 6345] = 175;
assign img[ 6346] = 172;
assign img[ 6347] = 172;
assign img[ 6348] = 174;
assign img[ 6349] = 174;
assign img[ 6350] = 175;
assign img[ 6351] = 174;
assign img[ 6352] = 192;
assign img[ 6353] = 176;
assign img[ 6354] = 175;
assign img[ 6355] = 172;
assign img[ 6356] = 174;
assign img[ 6357] = 172;
assign img[ 6358] = 175;
assign img[ 6359] = 176;
assign img[ 6360] = 175;
assign img[ 6361] = 176;
assign img[ 6362] = 192;
assign img[ 6363] = 172;
assign img[ 6364] = 172;
assign img[ 6365] = 180;
assign img[ 6366] = 175;
assign img[ 6367] = 169;
assign img[ 6368] = 177;
assign img[ 6369] = 180;
assign img[ 6370] = 173;
assign img[ 6371] = 184;
assign img[ 6372] = 174;
assign img[ 6373] = 175;
assign img[ 6374] = 172;
assign img[ 6375] = 175;
assign img[ 6376] = 174;
assign img[ 6377] = 172;
assign img[ 6378] = 176;
assign img[ 6379] = 174;
assign img[ 6380] = 175;
assign img[ 6381] = 172;
assign img[ 6382] = 174;
assign img[ 6383] = 167;
assign img[ 6384] = 175;
assign img[ 6385] = 173;
assign img[ 6386] = 175;
assign img[ 6387] = 174;
assign img[ 6388] = 164;
assign img[ 6389] = 173;
assign img[ 6390] = 175;
assign img[ 6391] = 175;
assign img[ 6392] = 172;
assign img[ 6393] = 172;
assign img[ 6394] = 174;
assign img[ 6395] = 175;
assign img[ 6396] = 176;
assign img[ 6397] = 174;
assign img[ 6398] = 174;
assign img[ 6399] = 171;
assign img[ 6400] = 175;
assign img[ 6401] = 196;
assign img[ 6402] = 192;
assign img[ 6403] = 194;
assign img[ 6404] = 198;
assign img[ 6405] = 192;
assign img[ 6406] = 192;
assign img[ 6407] = 198;
assign img[ 6408] = 197;
assign img[ 6409] = 207;
assign img[ 6410] = 206;
assign img[ 6411] = 216;
assign img[ 6412] = 208;
assign img[ 6413] = 208;
assign img[ 6414] = 204;
assign img[ 6415] = 208;
assign img[ 6416] = 208;
assign img[ 6417] = 208;
assign img[ 6418] = 208;
assign img[ 6419] = 207;
assign img[ 6420] = 215;
assign img[ 6421] = 207;
assign img[ 6422] = 222;
assign img[ 6423] = 208;
assign img[ 6424] = 208;
assign img[ 6425] = 208;
assign img[ 6426] = 208;
assign img[ 6427] = 207;
assign img[ 6428] = 208;
assign img[ 6429] = 208;
assign img[ 6430] = 208;
assign img[ 6431] = 208;
assign img[ 6432] = 207;
assign img[ 6433] = 208;
assign img[ 6434] = 208;
assign img[ 6435] = 207;
assign img[ 6436] = 208;
assign img[ 6437] = 206;
assign img[ 6438] = 208;
assign img[ 6439] = 208;
assign img[ 6440] = 207;
assign img[ 6441] = 208;
assign img[ 6442] = 199;
assign img[ 6443] = 204;
assign img[ 6444] = 196;
assign img[ 6445] = 192;
assign img[ 6446] = 192;
assign img[ 6447] = 192;
assign img[ 6448] = 192;
assign img[ 6449] = 192;
assign img[ 6450] = 194;
assign img[ 6451] = 192;
assign img[ 6452] = 194;
assign img[ 6453] = 192;
assign img[ 6454] = 176;
assign img[ 6455] = 192;
assign img[ 6456] = 192;
assign img[ 6457] = 192;
assign img[ 6458] = 193;
assign img[ 6459] = 181;
assign img[ 6460] = 176;
assign img[ 6461] = 181;
assign img[ 6462] = 192;
assign img[ 6463] = 176;
assign img[ 6464] = 192;
assign img[ 6465] = 176;
assign img[ 6466] = 181;
assign img[ 6467] = 176;
assign img[ 6468] = 173;
assign img[ 6469] = 175;
assign img[ 6470] = 179;
assign img[ 6471] = 173;
assign img[ 6472] = 173;
assign img[ 6473] = 192;
assign img[ 6474] = 179;
assign img[ 6475] = 193;
assign img[ 6476] = 183;
assign img[ 6477] = 176;
assign img[ 6478] = 180;
assign img[ 6479] = 192;
assign img[ 6480] = 175;
assign img[ 6481] = 175;
assign img[ 6482] = 175;
assign img[ 6483] = 181;
assign img[ 6484] = 192;
assign img[ 6485] = 192;
assign img[ 6486] = 192;
assign img[ 6487] = 175;
assign img[ 6488] = 175;
assign img[ 6489] = 192;
assign img[ 6490] = 176;
assign img[ 6491] = 192;
assign img[ 6492] = 173;
assign img[ 6493] = 172;
assign img[ 6494] = 175;
assign img[ 6495] = 172;
assign img[ 6496] = 172;
assign img[ 6497] = 174;
assign img[ 6498] = 192;
assign img[ 6499] = 172;
assign img[ 6500] = 174;
assign img[ 6501] = 172;
assign img[ 6502] = 192;
assign img[ 6503] = 174;
assign img[ 6504] = 180;
assign img[ 6505] = 170;
assign img[ 6506] = 172;
assign img[ 6507] = 172;
assign img[ 6508] = 173;
assign img[ 6509] = 172;
assign img[ 6510] = 173;
assign img[ 6511] = 175;
assign img[ 6512] = 172;
assign img[ 6513] = 174;
assign img[ 6514] = 177;
assign img[ 6515] = 172;
assign img[ 6516] = 173;
assign img[ 6517] = 166;
assign img[ 6518] = 176;
assign img[ 6519] = 169;
assign img[ 6520] = 172;
assign img[ 6521] = 168;
assign img[ 6522] = 169;
assign img[ 6523] = 170;
assign img[ 6524] = 175;
assign img[ 6525] = 168;
assign img[ 6526] = 174;
assign img[ 6527] = 173;
assign img[ 6528] = 176;
assign img[ 6529] = 172;
assign img[ 6530] = 169;
assign img[ 6531] = 165;
assign img[ 6532] = 177;
assign img[ 6533] = 169;
assign img[ 6534] = 177;
assign img[ 6535] = 178;
assign img[ 6536] = 172;
assign img[ 6537] = 192;
assign img[ 6538] = 194;
assign img[ 6539] = 194;
assign img[ 6540] = 194;
assign img[ 6541] = 194;
assign img[ 6542] = 199;
assign img[ 6543] = 200;
assign img[ 6544] = 196;
assign img[ 6545] = 198;
assign img[ 6546] = 194;
assign img[ 6547] = 197;
assign img[ 6548] = 199;
assign img[ 6549] = 198;
assign img[ 6550] = 199;
assign img[ 6551] = 195;
assign img[ 6552] = 198;
assign img[ 6553] = 199;
assign img[ 6554] = 200;
assign img[ 6555] = 194;
assign img[ 6556] = 198;
assign img[ 6557] = 194;
assign img[ 6558] = 194;
assign img[ 6559] = 194;
assign img[ 6560] = 198;
assign img[ 6561] = 195;
assign img[ 6562] = 194;
assign img[ 6563] = 199;
assign img[ 6564] = 198;
assign img[ 6565] = 198;
assign img[ 6566] = 198;
assign img[ 6567] = 198;
assign img[ 6568] = 194;
assign img[ 6569] = 196;
assign img[ 6570] = 192;
assign img[ 6571] = 194;
assign img[ 6572] = 176;
assign img[ 6573] = 192;
assign img[ 6574] = 166;
assign img[ 6575] = 167;
assign img[ 6576] = 175;
assign img[ 6577] = 167;
assign img[ 6578] = 167;
assign img[ 6579] = 168;
assign img[ 6580] = 162;
assign img[ 6581] = 164;
assign img[ 6582] = 167;
assign img[ 6583] = 166;
assign img[ 6584] = 168;
assign img[ 6585] = 167;
assign img[ 6586] = 167;
assign img[ 6587] = 168;
assign img[ 6588] = 164;
assign img[ 6589] = 164;
assign img[ 6590] = 154;
assign img[ 6591] = 172;
assign img[ 6592] = 161;
assign img[ 6593] = 165;
assign img[ 6594] = 161;
assign img[ 6595] = 160;
assign img[ 6596] = 161;
assign img[ 6597] = 164;
assign img[ 6598] = 164;
assign img[ 6599] = 151;
assign img[ 6600] = 158;
assign img[ 6601] = 161;
assign img[ 6602] = 160;
assign img[ 6603] = 161;
assign img[ 6604] = 162;
assign img[ 6605] = 165;
assign img[ 6606] = 161;
assign img[ 6607] = 168;
assign img[ 6608] = 161;
assign img[ 6609] = 160;
assign img[ 6610] = 164;
assign img[ 6611] = 162;
assign img[ 6612] = 161;
assign img[ 6613] = 164;
assign img[ 6614] = 156;
assign img[ 6615] = 162;
assign img[ 6616] = 156;
assign img[ 6617] = 163;
assign img[ 6618] = 160;
assign img[ 6619] = 158;
assign img[ 6620] = 159;
assign img[ 6621] = 157;
assign img[ 6622] = 162;
assign img[ 6623] = 160;
assign img[ 6624] = 164;
assign img[ 6625] = 158;
assign img[ 6626] = 154;
assign img[ 6627] = 160;
assign img[ 6628] = 168;
assign img[ 6629] = 153;
assign img[ 6630] = 147;
assign img[ 6631] = 165;
assign img[ 6632] = 158;
assign img[ 6633] = 162;
assign img[ 6634] = 168;
assign img[ 6635] = 144;
assign img[ 6636] = 159;
assign img[ 6637] = 160;
assign img[ 6638] = 161;
assign img[ 6639] = 161;
assign img[ 6640] = 154;
assign img[ 6641] = 153;
assign img[ 6642] = 162;
assign img[ 6643] = 164;
assign img[ 6644] = 148;
assign img[ 6645] = 156;
assign img[ 6646] = 154;
assign img[ 6647] = 146;
assign img[ 6648] = 144;
assign img[ 6649] = 156;
assign img[ 6650] = 160;
assign img[ 6651] = 154;
assign img[ 6652] = 161;
assign img[ 6653] = 152;
assign img[ 6654] = 146;
assign img[ 6655] = 162;
assign img[ 6656] = 155;
assign img[ 6657] = 166;
assign img[ 6658] = 170;
assign img[ 6659] = 162;
assign img[ 6660] = 160;
assign img[ 6661] = 151;
assign img[ 6662] = 164;
assign img[ 6663] = 165;
assign img[ 6664] = 169;
assign img[ 6665] = 174;
assign img[ 6666] = 175;
assign img[ 6667] = 177;
assign img[ 6668] = 174;
assign img[ 6669] = 174;
assign img[ 6670] = 182;
assign img[ 6671] = 176;
assign img[ 6672] = 176;
assign img[ 6673] = 192;
assign img[ 6674] = 168;
assign img[ 6675] = 176;
assign img[ 6676] = 175;
assign img[ 6677] = 192;
assign img[ 6678] = 182;
assign img[ 6679] = 176;
assign img[ 6680] = 175;
assign img[ 6681] = 192;
assign img[ 6682] = 176;
assign img[ 6683] = 180;
assign img[ 6684] = 192;
assign img[ 6685] = 182;
assign img[ 6686] = 174;
assign img[ 6687] = 176;
assign img[ 6688] = 192;
assign img[ 6689] = 192;
assign img[ 6690] = 192;
assign img[ 6691] = 176;
assign img[ 6692] = 178;
assign img[ 6693] = 174;
assign img[ 6694] = 180;
assign img[ 6695] = 174;
assign img[ 6696] = 176;
assign img[ 6697] = 192;
assign img[ 6698] = 175;
assign img[ 6699] = 172;
assign img[ 6700] = 168;
assign img[ 6701] = 166;
assign img[ 6702] = 151;
assign img[ 6703] = 151;
assign img[ 6704] = 152;
assign img[ 6705] = 151;
assign img[ 6706] = 144;
assign img[ 6707] = 151;
assign img[ 6708] = 151;
assign img[ 6709] = 152;
assign img[ 6710] = 160;
assign img[ 6711] = 144;
assign img[ 6712] = 152;
assign img[ 6713] = 160;
assign img[ 6714] = 158;
assign img[ 6715] = 151;
assign img[ 6716] = 152;
assign img[ 6717] = 143;
assign img[ 6718] = 160;
assign img[ 6719] = 141;
assign img[ 6720] = 144;
assign img[ 6721] = 143;
assign img[ 6722] = 140;
assign img[ 6723] = 144;
assign img[ 6724] = 144;
assign img[ 6725] = 148;
assign img[ 6726] = 144;
assign img[ 6727] = 145;
assign img[ 6728] = 148;
assign img[ 6729] = 142;
assign img[ 6730] = 144;
assign img[ 6731] = 149;
assign img[ 6732] = 152;
assign img[ 6733] = 137;
assign img[ 6734] = 146;
assign img[ 6735] = 145;
assign img[ 6736] = 144;
assign img[ 6737] = 150;
assign img[ 6738] = 144;
assign img[ 6739] = 144;
assign img[ 6740] = 150;
assign img[ 6741] = 153;
assign img[ 6742] = 149;
assign img[ 6743] = 144;
assign img[ 6744] = 153;
assign img[ 6745] = 154;
assign img[ 6746] = 142;
assign img[ 6747] = 146;
assign img[ 6748] = 149;
assign img[ 6749] = 145;
assign img[ 6750] = 148;
assign img[ 6751] = 149;
assign img[ 6752] = 141;
assign img[ 6753] = 143;
assign img[ 6754] = 140;
assign img[ 6755] = 144;
assign img[ 6756] = 147;
assign img[ 6757] = 144;
assign img[ 6758] = 141;
assign img[ 6759] = 144;
assign img[ 6760] = 149;
assign img[ 6761] = 143;
assign img[ 6762] = 142;
assign img[ 6763] = 142;
assign img[ 6764] = 143;
assign img[ 6765] = 144;
assign img[ 6766] = 152;
assign img[ 6767] = 141;
assign img[ 6768] = 141;
assign img[ 6769] = 135;
assign img[ 6770] = 144;
assign img[ 6771] = 140;
assign img[ 6772] = 144;
assign img[ 6773] = 148;
assign img[ 6774] = 139;
assign img[ 6775] = 140;
assign img[ 6776] = 148;
assign img[ 6777] = 137;
assign img[ 6778] = 148;
assign img[ 6779] = 141;
assign img[ 6780] = 144;
assign img[ 6781] = 143;
assign img[ 6782] = 142;
assign img[ 6783] = 140;
assign img[ 6784] = 143;
assign img[ 6785] = 180;
assign img[ 6786] = 173;
assign img[ 6787] = 172;
assign img[ 6788] = 171;
assign img[ 6789] = 175;
assign img[ 6790] = 172;
assign img[ 6791] = 168;
assign img[ 6792] = 174;
assign img[ 6793] = 192;
assign img[ 6794] = 194;
assign img[ 6795] = 194;
assign img[ 6796] = 194;
assign img[ 6797] = 192;
assign img[ 6798] = 192;
assign img[ 6799] = 198;
assign img[ 6800] = 192;
assign img[ 6801] = 194;
assign img[ 6802] = 194;
assign img[ 6803] = 198;
assign img[ 6804] = 194;
assign img[ 6805] = 192;
assign img[ 6806] = 194;
assign img[ 6807] = 192;
assign img[ 6808] = 192;
assign img[ 6809] = 195;
assign img[ 6810] = 192;
assign img[ 6811] = 198;
assign img[ 6812] = 193;
assign img[ 6813] = 194;
assign img[ 6814] = 194;
assign img[ 6815] = 194;
assign img[ 6816] = 192;
assign img[ 6817] = 198;
assign img[ 6818] = 195;
assign img[ 6819] = 192;
assign img[ 6820] = 194;
assign img[ 6821] = 194;
assign img[ 6822] = 198;
assign img[ 6823] = 194;
assign img[ 6824] = 194;
assign img[ 6825] = 194;
assign img[ 6826] = 195;
assign img[ 6827] = 192;
assign img[ 6828] = 183;
assign img[ 6829] = 192;
assign img[ 6830] = 192;
assign img[ 6831] = 168;
assign img[ 6832] = 167;
assign img[ 6833] = 164;
assign img[ 6834] = 168;
assign img[ 6835] = 168;
assign img[ 6836] = 162;
assign img[ 6837] = 163;
assign img[ 6838] = 168;
assign img[ 6839] = 166;
assign img[ 6840] = 163;
assign img[ 6841] = 160;
assign img[ 6842] = 165;
assign img[ 6843] = 167;
assign img[ 6844] = 164;
assign img[ 6845] = 166;
assign img[ 6846] = 162;
assign img[ 6847] = 148;
assign img[ 6848] = 154;
assign img[ 6849] = 153;
assign img[ 6850] = 155;
assign img[ 6851] = 158;
assign img[ 6852] = 153;
assign img[ 6853] = 154;
assign img[ 6854] = 168;
assign img[ 6855] = 156;
assign img[ 6856] = 160;
assign img[ 6857] = 148;
assign img[ 6858] = 160;
assign img[ 6859] = 155;
assign img[ 6860] = 156;
assign img[ 6861] = 153;
assign img[ 6862] = 156;
assign img[ 6863] = 156;
assign img[ 6864] = 156;
assign img[ 6865] = 159;
assign img[ 6866] = 156;
assign img[ 6867] = 161;
assign img[ 6868] = 152;
assign img[ 6869] = 157;
assign img[ 6870] = 152;
assign img[ 6871] = 152;
assign img[ 6872] = 153;
assign img[ 6873] = 152;
assign img[ 6874] = 161;
assign img[ 6875] = 156;
assign img[ 6876] = 156;
assign img[ 6877] = 153;
assign img[ 6878] = 157;
assign img[ 6879] = 153;
assign img[ 6880] = 161;
assign img[ 6881] = 156;
assign img[ 6882] = 153;
assign img[ 6883] = 156;
assign img[ 6884] = 155;
assign img[ 6885] = 160;
assign img[ 6886] = 162;
assign img[ 6887] = 153;
assign img[ 6888] = 153;
assign img[ 6889] = 154;
assign img[ 6890] = 157;
assign img[ 6891] = 157;
assign img[ 6892] = 156;
assign img[ 6893] = 156;
assign img[ 6894] = 152;
assign img[ 6895] = 154;
assign img[ 6896] = 157;
assign img[ 6897] = 153;
assign img[ 6898] = 156;
assign img[ 6899] = 161;
assign img[ 6900] = 156;
assign img[ 6901] = 143;
assign img[ 6902] = 149;
assign img[ 6903] = 148;
assign img[ 6904] = 156;
assign img[ 6905] = 150;
assign img[ 6906] = 151;
assign img[ 6907] = 157;
assign img[ 6908] = 150;
assign img[ 6909] = 153;
assign img[ 6910] = 149;
assign img[ 6911] = 151;
assign img[ 6912] = 150;
assign img[ 6913] = 160;
assign img[ 6914] = 164;
assign img[ 6915] = 159;
assign img[ 6916] = 160;
assign img[ 6917] = 163;
assign img[ 6918] = 160;
assign img[ 6919] = 156;
assign img[ 6920] = 160;
assign img[ 6921] = 170;
assign img[ 6922] = 180;
assign img[ 6923] = 176;
assign img[ 6924] = 176;
assign img[ 6925] = 192;
assign img[ 6926] = 192;
assign img[ 6927] = 180;
assign img[ 6928] = 176;
assign img[ 6929] = 192;
assign img[ 6930] = 180;
assign img[ 6931] = 192;
assign img[ 6932] = 192;
assign img[ 6933] = 174;
assign img[ 6934] = 192;
assign img[ 6935] = 179;
assign img[ 6936] = 192;
assign img[ 6937] = 173;
assign img[ 6938] = 180;
assign img[ 6939] = 179;
assign img[ 6940] = 192;
assign img[ 6941] = 173;
assign img[ 6942] = 192;
assign img[ 6943] = 192;
assign img[ 6944] = 192;
assign img[ 6945] = 172;
assign img[ 6946] = 192;
assign img[ 6947] = 176;
assign img[ 6948] = 177;
assign img[ 6949] = 180;
assign img[ 6950] = 176;
assign img[ 6951] = 177;
assign img[ 6952] = 177;
assign img[ 6953] = 178;
assign img[ 6954] = 192;
assign img[ 6955] = 176;
assign img[ 6956] = 177;
assign img[ 6957] = 172;
assign img[ 6958] = 165;
assign img[ 6959] = 160;
assign img[ 6960] = 150;
assign img[ 6961] = 155;
assign img[ 6962] = 152;
assign img[ 6963] = 153;
assign img[ 6964] = 161;
assign img[ 6965] = 152;
assign img[ 6966] = 154;
assign img[ 6967] = 145;
assign img[ 6968] = 150;
assign img[ 6969] = 160;
assign img[ 6970] = 140;
assign img[ 6971] = 152;
assign img[ 6972] = 148;
assign img[ 6973] = 146;
assign img[ 6974] = 150;
assign img[ 6975] = 152;
assign img[ 6976] = 153;
assign img[ 6977] = 153;
assign img[ 6978] = 147;
assign img[ 6979] = 148;
assign img[ 6980] = 148;
assign img[ 6981] = 153;
assign img[ 6982] = 149;
assign img[ 6983] = 152;
assign img[ 6984] = 153;
assign img[ 6985] = 148;
assign img[ 6986] = 154;
assign img[ 6987] = 148;
assign img[ 6988] = 144;
assign img[ 6989] = 145;
assign img[ 6990] = 156;
assign img[ 6991] = 143;
assign img[ 6992] = 145;
assign img[ 6993] = 144;
assign img[ 6994] = 144;
assign img[ 6995] = 149;
assign img[ 6996] = 160;
assign img[ 6997] = 142;
assign img[ 6998] = 145;
assign img[ 6999] = 148;
assign img[ 7000] = 142;
assign img[ 7001] = 149;
assign img[ 7002] = 141;
assign img[ 7003] = 145;
assign img[ 7004] = 151;
assign img[ 7005] = 141;
assign img[ 7006] = 141;
assign img[ 7007] = 143;
assign img[ 7008] = 145;
assign img[ 7009] = 149;
assign img[ 7010] = 156;
assign img[ 7011] = 144;
assign img[ 7012] = 149;
assign img[ 7013] = 143;
assign img[ 7014] = 149;
assign img[ 7015] = 143;
assign img[ 7016] = 141;
assign img[ 7017] = 148;
assign img[ 7018] = 143;
assign img[ 7019] = 150;
assign img[ 7020] = 153;
assign img[ 7021] = 145;
assign img[ 7022] = 142;
assign img[ 7023] = 144;
assign img[ 7024] = 140;
assign img[ 7025] = 137;
assign img[ 7026] = 150;
assign img[ 7027] = 148;
assign img[ 7028] = 148;
assign img[ 7029] = 140;
assign img[ 7030] = 148;
assign img[ 7031] = 144;
assign img[ 7032] = 142;
assign img[ 7033] = 149;
assign img[ 7034] = 141;
assign img[ 7035] = 144;
assign img[ 7036] = 142;
assign img[ 7037] = 142;
assign img[ 7038] = 143;
assign img[ 7039] = 144;
assign img[ 7040] = 144;
assign img[ 7041] = 147;
assign img[ 7042] = 157;
assign img[ 7043] = 153;
assign img[ 7044] = 148;
assign img[ 7045] = 154;
assign img[ 7046] = 157;
assign img[ 7047] = 153;
assign img[ 7048] = 148;
assign img[ 7049] = 165;
assign img[ 7050] = 173;
assign img[ 7051] = 166;
assign img[ 7052] = 165;
assign img[ 7053] = 165;
assign img[ 7054] = 170;
assign img[ 7055] = 169;
assign img[ 7056] = 165;
assign img[ 7057] = 167;
assign img[ 7058] = 177;
assign img[ 7059] = 173;
assign img[ 7060] = 168;
assign img[ 7061] = 166;
assign img[ 7062] = 181;
assign img[ 7063] = 173;
assign img[ 7064] = 173;
assign img[ 7065] = 173;
assign img[ 7066] = 173;
assign img[ 7067] = 169;
assign img[ 7068] = 162;
assign img[ 7069] = 169;
assign img[ 7070] = 165;
assign img[ 7071] = 172;
assign img[ 7072] = 167;
assign img[ 7073] = 167;
assign img[ 7074] = 173;
assign img[ 7075] = 164;
assign img[ 7076] = 169;
assign img[ 7077] = 173;
assign img[ 7078] = 169;
assign img[ 7079] = 169;
assign img[ 7080] = 166;
assign img[ 7081] = 169;
assign img[ 7082] = 170;
assign img[ 7083] = 169;
assign img[ 7084] = 161;
assign img[ 7085] = 173;
assign img[ 7086] = 172;
assign img[ 7087] = 165;
assign img[ 7088] = 141;
assign img[ 7089] = 145;
assign img[ 7090] = 144;
assign img[ 7091] = 153;
assign img[ 7092] = 143;
assign img[ 7093] = 141;
assign img[ 7094] = 140;
assign img[ 7095] = 137;
assign img[ 7096] = 149;
assign img[ 7097] = 137;
assign img[ 7098] = 143;
assign img[ 7099] = 145;
assign img[ 7100] = 137;
assign img[ 7101] = 143;
assign img[ 7102] = 145;
assign img[ 7103] = 141;
assign img[ 7104] = 137;
assign img[ 7105] = 149;
assign img[ 7106] = 141;
assign img[ 7107] = 141;
assign img[ 7108] = 133;
assign img[ 7109] = 141;
assign img[ 7110] = 141;
assign img[ 7111] = 145;
assign img[ 7112] = 145;
assign img[ 7113] = 140;
assign img[ 7114] = 143;
assign img[ 7115] = 137;
assign img[ 7116] = 137;
assign img[ 7117] = 145;
assign img[ 7118] = 138;
assign img[ 7119] = 141;
assign img[ 7120] = 137;
assign img[ 7121] = 140;
assign img[ 7122] = 136;
assign img[ 7123] = 148;
assign img[ 7124] = 141;
assign img[ 7125] = 136;
assign img[ 7126] = 137;
assign img[ 7127] = 136;
assign img[ 7128] = 144;
assign img[ 7129] = 136;
assign img[ 7130] = 140;
assign img[ 7131] = 140;
assign img[ 7132] = 140;
assign img[ 7133] = 140;
assign img[ 7134] = 141;
assign img[ 7135] = 137;
assign img[ 7136] = 138;
assign img[ 7137] = 142;
assign img[ 7138] = 137;
assign img[ 7139] = 133;
assign img[ 7140] = 140;
assign img[ 7141] = 136;
assign img[ 7142] = 136;
assign img[ 7143] = 140;
assign img[ 7144] = 132;
assign img[ 7145] = 138;
assign img[ 7146] = 137;
assign img[ 7147] = 133;
assign img[ 7148] = 132;
assign img[ 7149] = 133;
assign img[ 7150] = 137;
assign img[ 7151] = 142;
assign img[ 7152] = 136;
assign img[ 7153] = 132;
assign img[ 7154] = 137;
assign img[ 7155] = 136;
assign img[ 7156] = 136;
assign img[ 7157] = 132;
assign img[ 7158] = 132;
assign img[ 7159] = 136;
assign img[ 7160] = 140;
assign img[ 7161] = 136;
assign img[ 7162] = 132;
assign img[ 7163] = 136;
assign img[ 7164] = 132;
assign img[ 7165] = 142;
assign img[ 7166] = 140;
assign img[ 7167] = 133;
assign img[ 7168] = 133;
assign img[ 7169] = 156;
assign img[ 7170] = 156;
assign img[ 7171] = 146;
assign img[ 7172] = 156;
assign img[ 7173] = 152;
assign img[ 7174] = 150;
assign img[ 7175] = 147;
assign img[ 7176] = 160;
assign img[ 7177] = 162;
assign img[ 7178] = 168;
assign img[ 7179] = 172;
assign img[ 7180] = 166;
assign img[ 7181] = 171;
assign img[ 7182] = 175;
assign img[ 7183] = 177;
assign img[ 7184] = 161;
assign img[ 7185] = 165;
assign img[ 7186] = 172;
assign img[ 7187] = 170;
assign img[ 7188] = 173;
assign img[ 7189] = 172;
assign img[ 7190] = 170;
assign img[ 7191] = 169;
assign img[ 7192] = 170;
assign img[ 7193] = 177;
assign img[ 7194] = 166;
assign img[ 7195] = 172;
assign img[ 7196] = 167;
assign img[ 7197] = 165;
assign img[ 7198] = 162;
assign img[ 7199] = 176;
assign img[ 7200] = 163;
assign img[ 7201] = 165;
assign img[ 7202] = 166;
assign img[ 7203] = 182;
assign img[ 7204] = 172;
assign img[ 7205] = 169;
assign img[ 7206] = 170;
assign img[ 7207] = 169;
assign img[ 7208] = 169;
assign img[ 7209] = 168;
assign img[ 7210] = 164;
assign img[ 7211] = 168;
assign img[ 7212] = 169;
assign img[ 7213] = 164;
assign img[ 7214] = 164;
assign img[ 7215] = 162;
assign img[ 7216] = 153;
assign img[ 7217] = 144;
assign img[ 7218] = 151;
assign img[ 7219] = 141;
assign img[ 7220] = 145;
assign img[ 7221] = 149;
assign img[ 7222] = 145;
assign img[ 7223] = 140;
assign img[ 7224] = 144;
assign img[ 7225] = 141;
assign img[ 7226] = 140;
assign img[ 7227] = 146;
assign img[ 7228] = 141;
assign img[ 7229] = 145;
assign img[ 7230] = 144;
assign img[ 7231] = 143;
assign img[ 7232] = 148;
assign img[ 7233] = 145;
assign img[ 7234] = 138;
assign img[ 7235] = 146;
assign img[ 7236] = 145;
assign img[ 7237] = 146;
assign img[ 7238] = 143;
assign img[ 7239] = 140;
assign img[ 7240] = 140;
assign img[ 7241] = 143;
assign img[ 7242] = 148;
assign img[ 7243] = 136;
assign img[ 7244] = 143;
assign img[ 7245] = 142;
assign img[ 7246] = 134;
assign img[ 7247] = 144;
assign img[ 7248] = 144;
assign img[ 7249] = 145;
assign img[ 7250] = 138;
assign img[ 7251] = 141;
assign img[ 7252] = 133;
assign img[ 7253] = 143;
assign img[ 7254] = 135;
assign img[ 7255] = 133;
assign img[ 7256] = 135;
assign img[ 7257] = 138;
assign img[ 7258] = 140;
assign img[ 7259] = 134;
assign img[ 7260] = 133;
assign img[ 7261] = 135;
assign img[ 7262] = 136;
assign img[ 7263] = 134;
assign img[ 7264] = 136;
assign img[ 7265] = 140;
assign img[ 7266] = 140;
assign img[ 7267] = 141;
assign img[ 7268] = 140;
assign img[ 7269] = 141;
assign img[ 7270] = 137;
assign img[ 7271] = 141;
assign img[ 7272] = 134;
assign img[ 7273] = 140;
assign img[ 7274] = 141;
assign img[ 7275] = 133;
assign img[ 7276] = 133;
assign img[ 7277] = 142;
assign img[ 7278] = 146;
assign img[ 7279] = 135;
assign img[ 7280] = 136;
assign img[ 7281] = 137;
assign img[ 7282] = 133;
assign img[ 7283] = 134;
assign img[ 7284] = 133;
assign img[ 7285] = 135;
assign img[ 7286] = 140;
assign img[ 7287] = 131;
assign img[ 7288] = 140;
assign img[ 7289] = 136;
assign img[ 7290] = 130;
assign img[ 7291] = 140;
assign img[ 7292] = 138;
assign img[ 7293] = 132;
assign img[ 7294] = 133;
assign img[ 7295] = 135;
assign img[ 7296] = 136;
assign img[ 7297] = 144;
assign img[ 7298] = 138;
assign img[ 7299] = 142;
assign img[ 7300] = 144;
assign img[ 7301] = 141;
assign img[ 7302] = 145;
assign img[ 7303] = 148;
assign img[ 7304] = 142;
assign img[ 7305] = 156;
assign img[ 7306] = 153;
assign img[ 7307] = 157;
assign img[ 7308] = 164;
assign img[ 7309] = 156;
assign img[ 7310] = 160;
assign img[ 7311] = 158;
assign img[ 7312] = 156;
assign img[ 7313] = 169;
assign img[ 7314] = 157;
assign img[ 7315] = 161;
assign img[ 7316] = 162;
assign img[ 7317] = 156;
assign img[ 7318] = 164;
assign img[ 7319] = 164;
assign img[ 7320] = 156;
assign img[ 7321] = 161;
assign img[ 7322] = 158;
assign img[ 7323] = 158;
assign img[ 7324] = 162;
assign img[ 7325] = 163;
assign img[ 7326] = 164;
assign img[ 7327] = 168;
assign img[ 7328] = 159;
assign img[ 7329] = 156;
assign img[ 7330] = 159;
assign img[ 7331] = 168;
assign img[ 7332] = 160;
assign img[ 7333] = 164;
assign img[ 7334] = 156;
assign img[ 7335] = 164;
assign img[ 7336] = 168;
assign img[ 7337] = 157;
assign img[ 7338] = 158;
assign img[ 7339] = 164;
assign img[ 7340] = 168;
assign img[ 7341] = 164;
assign img[ 7342] = 150;
assign img[ 7343] = 149;
assign img[ 7344] = 154;
assign img[ 7345] = 143;
assign img[ 7346] = 136;
assign img[ 7347] = 132;
assign img[ 7348] = 136;
assign img[ 7349] = 132;
assign img[ 7350] = 135;
assign img[ 7351] = 135;
assign img[ 7352] = 137;
assign img[ 7353] = 132;
assign img[ 7354] = 132;
assign img[ 7355] = 134;
assign img[ 7356] = 128;
assign img[ 7357] = 132;
assign img[ 7358] = 128;
assign img[ 7359] = 134;
assign img[ 7360] = 132;
assign img[ 7361] = 140;
assign img[ 7362] = 128;
assign img[ 7363] = 132;
assign img[ 7364] = 128;
assign img[ 7365] = 134;
assign img[ 7366] = 132;
assign img[ 7367] = 129;
assign img[ 7368] = 135;
assign img[ 7369] = 128;
assign img[ 7370] = 133;
assign img[ 7371] = 134;
assign img[ 7372] = 128;
assign img[ 7373] = 131;
assign img[ 7374] = 138;
assign img[ 7375] = 138;
assign img[ 7376] = 128;
assign img[ 7377] = 138;
assign img[ 7378] = 128;
assign img[ 7379] = 136;
assign img[ 7380] = 129;
assign img[ 7381] = 129;
assign img[ 7382] = 132;
assign img[ 7383] = 132;
assign img[ 7384] = 128;
assign img[ 7385] = 132;
assign img[ 7386] = 134;
assign img[ 7387] = 132;
assign img[ 7388] = 134;
assign img[ 7389] = 130;
assign img[ 7390] = 135;
assign img[ 7391] = 134;
assign img[ 7392] = 128;
assign img[ 7393] = 131;
assign img[ 7394] = 132;
assign img[ 7395] = 130;
assign img[ 7396] = 130;
assign img[ 7397] = 128;
assign img[ 7398] = 132;
assign img[ 7399] = 128;
assign img[ 7400] = 132;
assign img[ 7401] = 128;
assign img[ 7402] = 130;
assign img[ 7403] = 131;
assign img[ 7404] = 128;
assign img[ 7405] = 134;
assign img[ 7406] = 128;
assign img[ 7407] = 134;
assign img[ 7408] = 130;
assign img[ 7409] = 134;
assign img[ 7410] = 135;
assign img[ 7411] = 130;
assign img[ 7412] = 132;
assign img[ 7413] = 128;
assign img[ 7414] = 130;
assign img[ 7415] = 129;
assign img[ 7416] = 128;
assign img[ 7417] = 130;
assign img[ 7418] = 134;
assign img[ 7419] = 132;
assign img[ 7420] = 132;
assign img[ 7421] = 128;
assign img[ 7422] = 131;
assign img[ 7423] = 130;
assign img[ 7424] = 128;
assign img[ 7425] = 128;
assign img[ 7426] = 128;
assign img[ 7427] = 128;
assign img[ 7428] = 109;
assign img[ 7429] = 128;
assign img[ 7430] = 128;
assign img[ 7431] = 128;
assign img[ 7432] = 128;
assign img[ 7433] = 132;
assign img[ 7434] = 133;
assign img[ 7435] = 129;
assign img[ 7436] = 132;
assign img[ 7437] = 137;
assign img[ 7438] = 128;
assign img[ 7439] = 134;
assign img[ 7440] = 132;
assign img[ 7441] = 137;
assign img[ 7442] = 136;
assign img[ 7443] = 132;
assign img[ 7444] = 133;
assign img[ 7445] = 133;
assign img[ 7446] = 137;
assign img[ 7447] = 128;
assign img[ 7448] = 133;
assign img[ 7449] = 129;
assign img[ 7450] = 136;
assign img[ 7451] = 128;
assign img[ 7452] = 128;
assign img[ 7453] = 133;
assign img[ 7454] = 137;
assign img[ 7455] = 137;
assign img[ 7456] = 133;
assign img[ 7457] = 131;
assign img[ 7458] = 128;
assign img[ 7459] = 132;
assign img[ 7460] = 135;
assign img[ 7461] = 129;
assign img[ 7462] = 130;
assign img[ 7463] = 136;
assign img[ 7464] = 140;
assign img[ 7465] = 130;
assign img[ 7466] = 129;
assign img[ 7467] = 135;
assign img[ 7468] = 132;
assign img[ 7469] = 129;
assign img[ 7470] = 130;
assign img[ 7471] = 128;
assign img[ 7472] = 132;
assign img[ 7473] = 128;
assign img[ 7474] = 128;
assign img[ 7475] = 110;
assign img[ 7476] = 105;
assign img[ 7477] = 110;
assign img[ 7478] = 100;
assign img[ 7479] = 101;
assign img[ 7480] = 104;
assign img[ 7481] = 106;
assign img[ 7482] = 105;
assign img[ 7483] = 102;
assign img[ 7484] = 97;
assign img[ 7485] = 101;
assign img[ 7486] = 102;
assign img[ 7487] = 106;
assign img[ 7488] = 97;
assign img[ 7489] = 100;
assign img[ 7490] = 102;
assign img[ 7491] = 106;
assign img[ 7492] = 96;
assign img[ 7493] = 96;
assign img[ 7494] = 97;
assign img[ 7495] = 97;
assign img[ 7496] = 98;
assign img[ 7497] = 102;
assign img[ 7498] = 108;
assign img[ 7499] = 97;
assign img[ 7500] = 96;
assign img[ 7501] = 103;
assign img[ 7502] = 97;
assign img[ 7503] = 98;
assign img[ 7504] = 102;
assign img[ 7505] = 105;
assign img[ 7506] = 97;
assign img[ 7507] = 108;
assign img[ 7508] = 108;
assign img[ 7509] = 97;
assign img[ 7510] = 97;
assign img[ 7511] = 103;
assign img[ 7512] = 101;
assign img[ 7513] = 97;
assign img[ 7514] = 98;
assign img[ 7515] = 98;
assign img[ 7516] = 98;
assign img[ 7517] = 100;
assign img[ 7518] = 98;
assign img[ 7519] = 101;
assign img[ 7520] = 101;
assign img[ 7521] = 106;
assign img[ 7522] = 101;
assign img[ 7523] = 101;
assign img[ 7524] = 104;
assign img[ 7525] = 99;
assign img[ 7526] = 104;
assign img[ 7527] = 97;
assign img[ 7528] = 101;
assign img[ 7529] = 98;
assign img[ 7530] = 100;
assign img[ 7531] = 98;
assign img[ 7532] = 97;
assign img[ 7533] = 90;
assign img[ 7534] = 100;
assign img[ 7535] = 97;
assign img[ 7536] = 99;
assign img[ 7537] = 98;
assign img[ 7538] = 99;
assign img[ 7539] = 100;
assign img[ 7540] = 100;
assign img[ 7541] = 98;
assign img[ 7542] = 104;
assign img[ 7543] = 97;
assign img[ 7544] = 96;
assign img[ 7545] = 98;
assign img[ 7546] = 99;
assign img[ 7547] = 105;
assign img[ 7548] = 90;
assign img[ 7549] = 97;
assign img[ 7550] = 97;
assign img[ 7551] = 99;
assign img[ 7552] = 96;
assign img[ 7553] = 146;
assign img[ 7554] = 150;
assign img[ 7555] = 144;
assign img[ 7556] = 143;
assign img[ 7557] = 148;
assign img[ 7558] = 144;
assign img[ 7559] = 139;
assign img[ 7560] = 161;
assign img[ 7561] = 160;
assign img[ 7562] = 161;
assign img[ 7563] = 161;
assign img[ 7564] = 161;
assign img[ 7565] = 161;
assign img[ 7566] = 161;
assign img[ 7567] = 163;
assign img[ 7568] = 161;
assign img[ 7569] = 168;
assign img[ 7570] = 165;
assign img[ 7571] = 163;
assign img[ 7572] = 161;
assign img[ 7573] = 163;
assign img[ 7574] = 160;
assign img[ 7575] = 160;
assign img[ 7576] = 173;
assign img[ 7577] = 164;
assign img[ 7578] = 170;
assign img[ 7579] = 168;
assign img[ 7580] = 161;
assign img[ 7581] = 168;
assign img[ 7582] = 161;
assign img[ 7583] = 161;
assign img[ 7584] = 164;
assign img[ 7585] = 161;
assign img[ 7586] = 162;
assign img[ 7587] = 169;
assign img[ 7588] = 161;
assign img[ 7589] = 161;
assign img[ 7590] = 162;
assign img[ 7591] = 161;
assign img[ 7592] = 168;
assign img[ 7593] = 169;
assign img[ 7594] = 161;
assign img[ 7595] = 167;
assign img[ 7596] = 161;
assign img[ 7597] = 162;
assign img[ 7598] = 161;
assign img[ 7599] = 176;
assign img[ 7600] = 164;
assign img[ 7601] = 160;
assign img[ 7602] = 143;
assign img[ 7603] = 145;
assign img[ 7604] = 137;
assign img[ 7605] = 137;
assign img[ 7606] = 136;
assign img[ 7607] = 132;
assign img[ 7608] = 136;
assign img[ 7609] = 140;
assign img[ 7610] = 140;
assign img[ 7611] = 140;
assign img[ 7612] = 133;
assign img[ 7613] = 130;
assign img[ 7614] = 140;
assign img[ 7615] = 136;
assign img[ 7616] = 138;
assign img[ 7617] = 136;
assign img[ 7618] = 137;
assign img[ 7619] = 130;
assign img[ 7620] = 139;
assign img[ 7621] = 136;
assign img[ 7622] = 142;
assign img[ 7623] = 136;
assign img[ 7624] = 132;
assign img[ 7625] = 132;
assign img[ 7626] = 132;
assign img[ 7627] = 132;
assign img[ 7628] = 132;
assign img[ 7629] = 132;
assign img[ 7630] = 134;
assign img[ 7631] = 138;
assign img[ 7632] = 138;
assign img[ 7633] = 136;
assign img[ 7634] = 132;
assign img[ 7635] = 138;
assign img[ 7636] = 138;
assign img[ 7637] = 128;
assign img[ 7638] = 134;
assign img[ 7639] = 128;
assign img[ 7640] = 130;
assign img[ 7641] = 131;
assign img[ 7642] = 134;
assign img[ 7643] = 134;
assign img[ 7644] = 138;
assign img[ 7645] = 128;
assign img[ 7646] = 134;
assign img[ 7647] = 136;
assign img[ 7648] = 137;
assign img[ 7649] = 129;
assign img[ 7650] = 134;
assign img[ 7651] = 133;
assign img[ 7652] = 128;
assign img[ 7653] = 131;
assign img[ 7654] = 136;
assign img[ 7655] = 136;
assign img[ 7656] = 130;
assign img[ 7657] = 139;
assign img[ 7658] = 140;
assign img[ 7659] = 134;
assign img[ 7660] = 129;
assign img[ 7661] = 128;
assign img[ 7662] = 130;
assign img[ 7663] = 135;
assign img[ 7664] = 129;
assign img[ 7665] = 131;
assign img[ 7666] = 131;
assign img[ 7667] = 129;
assign img[ 7668] = 132;
assign img[ 7669] = 129;
assign img[ 7670] = 132;
assign img[ 7671] = 132;
assign img[ 7672] = 129;
assign img[ 7673] = 130;
assign img[ 7674] = 136;
assign img[ 7675] = 136;
assign img[ 7676] = 128;
assign img[ 7677] = 131;
assign img[ 7678] = 135;
assign img[ 7679] = 136;
assign img[ 7680] = 136;
assign img[ 7681] = 137;
assign img[ 7682] = 138;
assign img[ 7683] = 132;
assign img[ 7684] = 139;
assign img[ 7685] = 129;
assign img[ 7686] = 136;
assign img[ 7687] = 136;
assign img[ 7688] = 142;
assign img[ 7689] = 148;
assign img[ 7690] = 144;
assign img[ 7691] = 153;
assign img[ 7692] = 148;
assign img[ 7693] = 152;
assign img[ 7694] = 153;
assign img[ 7695] = 153;
assign img[ 7696] = 153;
assign img[ 7697] = 156;
assign img[ 7698] = 160;
assign img[ 7699] = 161;
assign img[ 7700] = 153;
assign img[ 7701] = 149;
assign img[ 7702] = 154;
assign img[ 7703] = 160;
assign img[ 7704] = 140;
assign img[ 7705] = 150;
assign img[ 7706] = 150;
assign img[ 7707] = 147;
assign img[ 7708] = 147;
assign img[ 7709] = 148;
assign img[ 7710] = 154;
assign img[ 7711] = 153;
assign img[ 7712] = 161;
assign img[ 7713] = 156;
assign img[ 7714] = 160;
assign img[ 7715] = 164;
assign img[ 7716] = 153;
assign img[ 7717] = 153;
assign img[ 7718] = 154;
assign img[ 7719] = 146;
assign img[ 7720] = 152;
assign img[ 7721] = 164;
assign img[ 7722] = 149;
assign img[ 7723] = 160;
assign img[ 7724] = 152;
assign img[ 7725] = 161;
assign img[ 7726] = 148;
assign img[ 7727] = 150;
assign img[ 7728] = 154;
assign img[ 7729] = 144;
assign img[ 7730] = 141;
assign img[ 7731] = 133;
assign img[ 7732] = 129;
assign img[ 7733] = 130;
assign img[ 7734] = 135;
assign img[ 7735] = 132;
assign img[ 7736] = 128;
assign img[ 7737] = 128;
assign img[ 7738] = 129;
assign img[ 7739] = 128;
assign img[ 7740] = 133;
assign img[ 7741] = 129;
assign img[ 7742] = 128;
assign img[ 7743] = 128;
assign img[ 7744] = 128;
assign img[ 7745] = 129;
assign img[ 7746] = 130;
assign img[ 7747] = 129;
assign img[ 7748] = 129;
assign img[ 7749] = 128;
assign img[ 7750] = 128;
assign img[ 7751] = 130;
assign img[ 7752] = 129;
assign img[ 7753] = 128;
assign img[ 7754] = 128;
assign img[ 7755] = 128;
assign img[ 7756] = 128;
assign img[ 7757] = 129;
assign img[ 7758] = 128;
assign img[ 7759] = 128;
assign img[ 7760] = 128;
assign img[ 7761] = 128;
assign img[ 7762] = 128;
assign img[ 7763] = 130;
assign img[ 7764] = 128;
assign img[ 7765] = 130;
assign img[ 7766] = 128;
assign img[ 7767] = 128;
assign img[ 7768] = 128;
assign img[ 7769] = 128;
assign img[ 7770] = 128;
assign img[ 7771] = 128;
assign img[ 7772] = 130;
assign img[ 7773] = 128;
assign img[ 7774] = 128;
assign img[ 7775] = 128;
assign img[ 7776] = 128;
assign img[ 7777] = 128;
assign img[ 7778] = 128;
assign img[ 7779] = 128;
assign img[ 7780] = 128;
assign img[ 7781] = 128;
assign img[ 7782] = 128;
assign img[ 7783] = 128;
assign img[ 7784] = 128;
assign img[ 7785] = 128;
assign img[ 7786] = 128;
assign img[ 7787] = 128;
assign img[ 7788] = 128;
assign img[ 7789] = 128;
assign img[ 7790] = 130;
assign img[ 7791] = 128;
assign img[ 7792] = 111;
assign img[ 7793] = 128;
assign img[ 7794] = 128;
assign img[ 7795] = 128;
assign img[ 7796] = 128;
assign img[ 7797] = 128;
assign img[ 7798] = 128;
assign img[ 7799] = 128;
assign img[ 7800] = 128;
assign img[ 7801] = 128;
assign img[ 7802] = 128;
assign img[ 7803] = 128;
assign img[ 7804] = 128;
assign img[ 7805] = 128;
assign img[ 7806] = 128;
assign img[ 7807] = 128;
assign img[ 7808] = 128;
assign img[ 7809] = 128;
assign img[ 7810] = 128;
assign img[ 7811] = 128;
assign img[ 7812] = 104;
assign img[ 7813] = 128;
assign img[ 7814] = 128;
assign img[ 7815] = 112;
assign img[ 7816] = 128;
assign img[ 7817] = 131;
assign img[ 7818] = 136;
assign img[ 7819] = 143;
assign img[ 7820] = 130;
assign img[ 7821] = 137;
assign img[ 7822] = 133;
assign img[ 7823] = 140;
assign img[ 7824] = 140;
assign img[ 7825] = 142;
assign img[ 7826] = 138;
assign img[ 7827] = 141;
assign img[ 7828] = 141;
assign img[ 7829] = 146;
assign img[ 7830] = 142;
assign img[ 7831] = 137;
assign img[ 7832] = 141;
assign img[ 7833] = 137;
assign img[ 7834] = 139;
assign img[ 7835] = 138;
assign img[ 7836] = 132;
assign img[ 7837] = 136;
assign img[ 7838] = 141;
assign img[ 7839] = 143;
assign img[ 7840] = 141;
assign img[ 7841] = 135;
assign img[ 7842] = 137;
assign img[ 7843] = 141;
assign img[ 7844] = 137;
assign img[ 7845] = 141;
assign img[ 7846] = 137;
assign img[ 7847] = 141;
assign img[ 7848] = 141;
assign img[ 7849] = 145;
assign img[ 7850] = 134;
assign img[ 7851] = 143;
assign img[ 7852] = 145;
assign img[ 7853] = 138;
assign img[ 7854] = 137;
assign img[ 7855] = 136;
assign img[ 7856] = 137;
assign img[ 7857] = 135;
assign img[ 7858] = 129;
assign img[ 7859] = 130;
assign img[ 7860] = 128;
assign img[ 7861] = 128;
assign img[ 7862] = 113;
assign img[ 7863] = 106;
assign img[ 7864] = 113;
assign img[ 7865] = 128;
assign img[ 7866] = 105;
assign img[ 7867] = 108;
assign img[ 7868] = 128;
assign img[ 7869] = 109;
assign img[ 7870] = 107;
assign img[ 7871] = 129;
assign img[ 7872] = 101;
assign img[ 7873] = 105;
assign img[ 7874] = 105;
assign img[ 7875] = 105;
assign img[ 7876] = 105;
assign img[ 7877] = 113;
assign img[ 7878] = 112;
assign img[ 7879] = 114;
assign img[ 7880] = 108;
assign img[ 7881] = 105;
assign img[ 7882] = 106;
assign img[ 7883] = 104;
assign img[ 7884] = 101;
assign img[ 7885] = 105;
assign img[ 7886] = 108;
assign img[ 7887] = 128;
assign img[ 7888] = 104;
assign img[ 7889] = 106;
assign img[ 7890] = 104;
assign img[ 7891] = 110;
assign img[ 7892] = 112;
assign img[ 7893] = 109;
assign img[ 7894] = 111;
assign img[ 7895] = 103;
assign img[ 7896] = 102;
assign img[ 7897] = 103;
assign img[ 7898] = 104;
assign img[ 7899] = 102;
assign img[ 7900] = 103;
assign img[ 7901] = 105;
assign img[ 7902] = 103;
assign img[ 7903] = 106;
assign img[ 7904] = 102;
assign img[ 7905] = 99;
assign img[ 7906] = 102;
assign img[ 7907] = 100;
assign img[ 7908] = 112;
assign img[ 7909] = 103;
assign img[ 7910] = 128;
assign img[ 7911] = 101;
assign img[ 7912] = 97;
assign img[ 7913] = 107;
assign img[ 7914] = 100;
assign img[ 7915] = 106;
assign img[ 7916] = 100;
assign img[ 7917] = 106;
assign img[ 7918] = 106;
assign img[ 7919] = 105;
assign img[ 7920] = 105;
assign img[ 7921] = 102;
assign img[ 7922] = 104;
assign img[ 7923] = 99;
assign img[ 7924] = 108;
assign img[ 7925] = 97;
assign img[ 7926] = 98;
assign img[ 7927] = 110;
assign img[ 7928] = 104;
assign img[ 7929] = 102;
assign img[ 7930] = 101;
assign img[ 7931] = 102;
assign img[ 7932] = 104;
assign img[ 7933] = 112;
assign img[ 7934] = 100;
assign img[ 7935] = 99;
assign img[ 7936] = 108;
assign img[ 7937] = 144;
assign img[ 7938] = 147;
assign img[ 7939] = 140;
assign img[ 7940] = 150;
assign img[ 7941] = 144;
assign img[ 7942] = 142;
assign img[ 7943] = 148;
assign img[ 7944] = 143;
assign img[ 7945] = 142;
assign img[ 7946] = 161;
assign img[ 7947] = 162;
assign img[ 7948] = 161;
assign img[ 7949] = 149;
assign img[ 7950] = 161;
assign img[ 7951] = 167;
assign img[ 7952] = 161;
assign img[ 7953] = 162;
assign img[ 7954] = 164;
assign img[ 7955] = 161;
assign img[ 7956] = 162;
assign img[ 7957] = 164;
assign img[ 7958] = 161;
assign img[ 7959] = 164;
assign img[ 7960] = 165;
assign img[ 7961] = 153;
assign img[ 7962] = 156;
assign img[ 7963] = 161;
assign img[ 7964] = 161;
assign img[ 7965] = 165;
assign img[ 7966] = 157;
assign img[ 7967] = 164;
assign img[ 7968] = 160;
assign img[ 7969] = 153;
assign img[ 7970] = 160;
assign img[ 7971] = 153;
assign img[ 7972] = 164;
assign img[ 7973] = 160;
assign img[ 7974] = 161;
assign img[ 7975] = 164;
assign img[ 7976] = 162;
assign img[ 7977] = 162;
assign img[ 7978] = 165;
assign img[ 7979] = 170;
assign img[ 7980] = 165;
assign img[ 7981] = 161;
assign img[ 7982] = 162;
assign img[ 7983] = 165;
assign img[ 7984] = 157;
assign img[ 7985] = 160;
assign img[ 7986] = 153;
assign img[ 7987] = 165;
assign img[ 7988] = 153;
assign img[ 7989] = 149;
assign img[ 7990] = 142;
assign img[ 7991] = 137;
assign img[ 7992] = 132;
assign img[ 7993] = 129;
assign img[ 7994] = 133;
assign img[ 7995] = 136;
assign img[ 7996] = 141;
assign img[ 7997] = 137;
assign img[ 7998] = 129;
assign img[ 7999] = 133;
assign img[ 8000] = 129;
assign img[ 8001] = 133;
assign img[ 8002] = 129;
assign img[ 8003] = 137;
assign img[ 8004] = 128;
assign img[ 8005] = 141;
assign img[ 8006] = 132;
assign img[ 8007] = 129;
assign img[ 8008] = 133;
assign img[ 8009] = 133;
assign img[ 8010] = 129;
assign img[ 8011] = 130;
assign img[ 8012] = 132;
assign img[ 8013] = 130;
assign img[ 8014] = 132;
assign img[ 8015] = 130;
assign img[ 8016] = 128;
assign img[ 8017] = 128;
assign img[ 8018] = 131;
assign img[ 8019] = 134;
assign img[ 8020] = 129;
assign img[ 8021] = 128;
assign img[ 8022] = 132;
assign img[ 8023] = 128;
assign img[ 8024] = 128;
assign img[ 8025] = 134;
assign img[ 8026] = 128;
assign img[ 8027] = 128;
assign img[ 8028] = 134;
assign img[ 8029] = 132;
assign img[ 8030] = 128;
assign img[ 8031] = 128;
assign img[ 8032] = 128;
assign img[ 8033] = 135;
assign img[ 8034] = 137;
assign img[ 8035] = 128;
assign img[ 8036] = 128;
assign img[ 8037] = 132;
assign img[ 8038] = 128;
assign img[ 8039] = 128;
assign img[ 8040] = 128;
assign img[ 8041] = 128;
assign img[ 8042] = 130;
assign img[ 8043] = 135;
assign img[ 8044] = 128;
assign img[ 8045] = 132;
assign img[ 8046] = 132;
assign img[ 8047] = 133;
assign img[ 8048] = 128;
assign img[ 8049] = 128;
assign img[ 8050] = 132;
assign img[ 8051] = 128;
assign img[ 8052] = 132;
assign img[ 8053] = 128;
assign img[ 8054] = 132;
assign img[ 8055] = 132;
assign img[ 8056] = 128;
assign img[ 8057] = 128;
assign img[ 8058] = 128;
assign img[ 8059] = 128;
assign img[ 8060] = 128;
assign img[ 8061] = 128;
assign img[ 8062] = 128;
assign img[ 8063] = 128;
assign img[ 8064] = 129;
assign img[ 8065] = 148;
assign img[ 8066] = 144;
assign img[ 8067] = 148;
assign img[ 8068] = 153;
assign img[ 8069] = 144;
assign img[ 8070] = 152;
assign img[ 8071] = 160;
assign img[ 8072] = 150;
assign img[ 8073] = 161;
assign img[ 8074] = 165;
assign img[ 8075] = 164;
assign img[ 8076] = 162;
assign img[ 8077] = 164;
assign img[ 8078] = 169;
assign img[ 8079] = 169;
assign img[ 8080] = 161;
assign img[ 8081] = 169;
assign img[ 8082] = 173;
assign img[ 8083] = 163;
assign img[ 8084] = 175;
assign img[ 8085] = 165;
assign img[ 8086] = 169;
assign img[ 8087] = 162;
assign img[ 8088] = 161;
assign img[ 8089] = 164;
assign img[ 8090] = 171;
assign img[ 8091] = 169;
assign img[ 8092] = 173;
assign img[ 8093] = 169;
assign img[ 8094] = 168;
assign img[ 8095] = 164;
assign img[ 8096] = 169;
assign img[ 8097] = 169;
assign img[ 8098] = 165;
assign img[ 8099] = 173;
assign img[ 8100] = 162;
assign img[ 8101] = 169;
assign img[ 8102] = 169;
assign img[ 8103] = 171;
assign img[ 8104] = 169;
assign img[ 8105] = 169;
assign img[ 8106] = 171;
assign img[ 8107] = 169;
assign img[ 8108] = 168;
assign img[ 8109] = 173;
assign img[ 8110] = 165;
assign img[ 8111] = 169;
assign img[ 8112] = 169;
assign img[ 8113] = 168;
assign img[ 8114] = 172;
assign img[ 8115] = 162;
assign img[ 8116] = 165;
assign img[ 8117] = 161;
assign img[ 8118] = 161;
assign img[ 8119] = 153;
assign img[ 8120] = 139;
assign img[ 8121] = 143;
assign img[ 8122] = 139;
assign img[ 8123] = 145;
assign img[ 8124] = 144;
assign img[ 8125] = 145;
assign img[ 8126] = 144;
assign img[ 8127] = 138;
assign img[ 8128] = 137;
assign img[ 8129] = 138;
assign img[ 8130] = 141;
assign img[ 8131] = 146;
assign img[ 8132] = 139;
assign img[ 8133] = 145;
assign img[ 8134] = 141;
assign img[ 8135] = 145;
assign img[ 8136] = 137;
assign img[ 8137] = 135;
assign img[ 8138] = 141;
assign img[ 8139] = 145;
assign img[ 8140] = 136;
assign img[ 8141] = 143;
assign img[ 8142] = 148;
assign img[ 8143] = 137;
assign img[ 8144] = 139;
assign img[ 8145] = 141;
assign img[ 8146] = 137;
assign img[ 8147] = 138;
assign img[ 8148] = 146;
assign img[ 8149] = 140;
assign img[ 8150] = 140;
assign img[ 8151] = 137;
assign img[ 8152] = 133;
assign img[ 8153] = 141;
assign img[ 8154] = 143;
assign img[ 8155] = 140;
assign img[ 8156] = 139;
assign img[ 8157] = 137;
assign img[ 8158] = 140;
assign img[ 8159] = 140;
assign img[ 8160] = 131;
assign img[ 8161] = 137;
assign img[ 8162] = 141;
assign img[ 8163] = 140;
assign img[ 8164] = 139;
assign img[ 8165] = 145;
assign img[ 8166] = 134;
assign img[ 8167] = 139;
assign img[ 8168] = 137;
assign img[ 8169] = 141;
assign img[ 8170] = 137;
assign img[ 8171] = 141;
assign img[ 8172] = 139;
assign img[ 8173] = 141;
assign img[ 8174] = 137;
assign img[ 8175] = 140;
assign img[ 8176] = 137;
assign img[ 8177] = 131;
assign img[ 8178] = 138;
assign img[ 8179] = 137;
assign img[ 8180] = 129;
assign img[ 8181] = 133;
assign img[ 8182] = 139;
assign img[ 8183] = 137;
assign img[ 8184] = 135;
assign img[ 8185] = 129;
assign img[ 8186] = 140;
assign img[ 8187] = 136;
assign img[ 8188] = 145;
assign img[ 8189] = 135;
assign img[ 8190] = 140;
assign img[ 8191] = 137;
assign img[ 8192] = 53;
assign img[ 8193] = 89;
assign img[ 8194] = 84;
assign img[ 8195] = 80;
assign img[ 8196] = 87;
assign img[ 8197] = 86;
assign img[ 8198] = 88;
assign img[ 8199] = 80;
assign img[ 8200] = 92;
assign img[ 8201] = 88;
assign img[ 8202] = 103;
assign img[ 8203] = 104;
assign img[ 8204] = 101;
assign img[ 8205] = 104;
assign img[ 8206] = 99;
assign img[ 8207] = 104;
assign img[ 8208] = 108;
assign img[ 8209] = 104;
assign img[ 8210] = 107;
assign img[ 8211] = 103;
assign img[ 8212] = 104;
assign img[ 8213] = 104;
assign img[ 8214] = 108;
assign img[ 8215] = 105;
assign img[ 8216] = 103;
assign img[ 8217] = 101;
assign img[ 8218] = 110;
assign img[ 8219] = 104;
assign img[ 8220] = 101;
assign img[ 8221] = 106;
assign img[ 8222] = 104;
assign img[ 8223] = 107;
assign img[ 8224] = 104;
assign img[ 8225] = 105;
assign img[ 8226] = 102;
assign img[ 8227] = 128;
assign img[ 8228] = 104;
assign img[ 8229] = 103;
assign img[ 8230] = 103;
assign img[ 8231] = 101;
assign img[ 8232] = 103;
assign img[ 8233] = 100;
assign img[ 8234] = 103;
assign img[ 8235] = 107;
assign img[ 8236] = 102;
assign img[ 8237] = 105;
assign img[ 8238] = 101;
assign img[ 8239] = 110;
assign img[ 8240] = 110;
assign img[ 8241] = 128;
assign img[ 8242] = 103;
assign img[ 8243] = 103;
assign img[ 8244] = 102;
assign img[ 8245] = 97;
assign img[ 8246] = 108;
assign img[ 8247] = 98;
assign img[ 8248] = 99;
assign img[ 8249] = 96;
assign img[ 8250] = 86;
assign img[ 8251] = 79;
assign img[ 8252] = 85;
assign img[ 8253] = 80;
assign img[ 8254] = 86;
assign img[ 8255] = 80;
assign img[ 8256] = 78;
assign img[ 8257] = 78;
assign img[ 8258] = 74;
assign img[ 8259] = 79;
assign img[ 8260] = 76;
assign img[ 8261] = 77;
assign img[ 8262] = 75;
assign img[ 8263] = 83;
assign img[ 8264] = 85;
assign img[ 8265] = 77;
assign img[ 8266] = 79;
assign img[ 8267] = 78;
assign img[ 8268] = 74;
assign img[ 8269] = 76;
assign img[ 8270] = 77;
assign img[ 8271] = 78;
assign img[ 8272] = 78;
assign img[ 8273] = 74;
assign img[ 8274] = 70;
assign img[ 8275] = 79;
assign img[ 8276] = 76;
assign img[ 8277] = 78;
assign img[ 8278] = 80;
assign img[ 8279] = 76;
assign img[ 8280] = 76;
assign img[ 8281] = 84;
assign img[ 8282] = 77;
assign img[ 8283] = 78;
assign img[ 8284] = 71;
assign img[ 8285] = 76;
assign img[ 8286] = 70;
assign img[ 8287] = 68;
assign img[ 8288] = 68;
assign img[ 8289] = 70;
assign img[ 8290] = 70;
assign img[ 8291] = 76;
assign img[ 8292] = 70;
assign img[ 8293] = 70;
assign img[ 8294] = 72;
assign img[ 8295] = 72;
assign img[ 8296] = 78;
assign img[ 8297] = 76;
assign img[ 8298] = 72;
assign img[ 8299] = 68;
assign img[ 8300] = 68;
assign img[ 8301] = 70;
assign img[ 8302] = 68;
assign img[ 8303] = 76;
assign img[ 8304] = 70;
assign img[ 8305] = 74;
assign img[ 8306] = 71;
assign img[ 8307] = 72;
assign img[ 8308] = 68;
assign img[ 8309] = 76;
assign img[ 8310] = 72;
assign img[ 8311] = 68;
assign img[ 8312] = 69;
assign img[ 8313] = 70;
assign img[ 8314] = 70;
assign img[ 8315] = 68;
assign img[ 8316] = 76;
assign img[ 8317] = 68;
assign img[ 8318] = 71;
assign img[ 8319] = 71;
assign img[ 8320] = 76;
assign img[ 8321] = 102;
assign img[ 8322] = 100;
assign img[ 8323] = 96;
assign img[ 8324] = 94;
assign img[ 8325] = 101;
assign img[ 8326] = 98;
assign img[ 8327] = 98;
assign img[ 8328] = 105;
assign img[ 8329] = 104;
assign img[ 8330] = 104;
assign img[ 8331] = 128;
assign img[ 8332] = 128;
assign img[ 8333] = 128;
assign img[ 8334] = 110;
assign img[ 8335] = 128;
assign img[ 8336] = 128;
assign img[ 8337] = 128;
assign img[ 8338] = 128;
assign img[ 8339] = 128;
assign img[ 8340] = 112;
assign img[ 8341] = 128;
assign img[ 8342] = 128;
assign img[ 8343] = 112;
assign img[ 8344] = 128;
assign img[ 8345] = 128;
assign img[ 8346] = 128;
assign img[ 8347] = 128;
assign img[ 8348] = 128;
assign img[ 8349] = 128;
assign img[ 8350] = 128;
assign img[ 8351] = 128;
assign img[ 8352] = 128;
assign img[ 8353] = 128;
assign img[ 8354] = 128;
assign img[ 8355] = 128;
assign img[ 8356] = 108;
assign img[ 8357] = 128;
assign img[ 8358] = 128;
assign img[ 8359] = 128;
assign img[ 8360] = 128;
assign img[ 8361] = 130;
assign img[ 8362] = 128;
assign img[ 8363] = 128;
assign img[ 8364] = 128;
assign img[ 8365] = 128;
assign img[ 8366] = 128;
assign img[ 8367] = 128;
assign img[ 8368] = 128;
assign img[ 8369] = 128;
assign img[ 8370] = 128;
assign img[ 8371] = 128;
assign img[ 8372] = 128;
assign img[ 8373] = 128;
assign img[ 8374] = 128;
assign img[ 8375] = 112;
assign img[ 8376] = 110;
assign img[ 8377] = 102;
assign img[ 8378] = 96;
assign img[ 8379] = 96;
assign img[ 8380] = 92;
assign img[ 8381] = 90;
assign img[ 8382] = 89;
assign img[ 8383] = 96;
assign img[ 8384] = 86;
assign img[ 8385] = 97;
assign img[ 8386] = 84;
assign img[ 8387] = 86;
assign img[ 8388] = 87;
assign img[ 8389] = 84;
assign img[ 8390] = 97;
assign img[ 8391] = 84;
assign img[ 8392] = 91;
assign img[ 8393] = 92;
assign img[ 8394] = 84;
assign img[ 8395] = 93;
assign img[ 8396] = 94;
assign img[ 8397] = 86;
assign img[ 8398] = 86;
assign img[ 8399] = 86;
assign img[ 8400] = 96;
assign img[ 8401] = 88;
assign img[ 8402] = 92;
assign img[ 8403] = 86;
assign img[ 8404] = 94;
assign img[ 8405] = 86;
assign img[ 8406] = 80;
assign img[ 8407] = 94;
assign img[ 8408] = 94;
assign img[ 8409] = 92;
assign img[ 8410] = 92;
assign img[ 8411] = 85;
assign img[ 8412] = 84;
assign img[ 8413] = 88;
assign img[ 8414] = 96;
assign img[ 8415] = 88;
assign img[ 8416] = 84;
assign img[ 8417] = 84;
assign img[ 8418] = 88;
assign img[ 8419] = 95;
assign img[ 8420] = 87;
assign img[ 8421] = 88;
assign img[ 8422] = 86;
assign img[ 8423] = 88;
assign img[ 8424] = 92;
assign img[ 8425] = 86;
assign img[ 8426] = 84;
assign img[ 8427] = 92;
assign img[ 8428] = 91;
assign img[ 8429] = 90;
assign img[ 8430] = 84;
assign img[ 8431] = 92;
assign img[ 8432] = 92;
assign img[ 8433] = 85;
assign img[ 8434] = 84;
assign img[ 8435] = 84;
assign img[ 8436] = 84;
assign img[ 8437] = 85;
assign img[ 8438] = 84;
assign img[ 8439] = 92;
assign img[ 8440] = 88;
assign img[ 8441] = 84;
assign img[ 8442] = 84;
assign img[ 8443] = 84;
assign img[ 8444] = 80;
assign img[ 8445] = 87;
assign img[ 8446] = 96;
assign img[ 8447] = 83;
assign img[ 8448] = 84;
assign img[ 8449] = 102;
assign img[ 8450] = 108;
assign img[ 8451] = 104;
assign img[ 8452] = 102;
assign img[ 8453] = 102;
assign img[ 8454] = 108;
assign img[ 8455] = 110;
assign img[ 8456] = 128;
assign img[ 8457] = 110;
assign img[ 8458] = 130;
assign img[ 8459] = 128;
assign img[ 8460] = 132;
assign img[ 8461] = 130;
assign img[ 8462] = 128;
assign img[ 8463] = 134;
assign img[ 8464] = 132;
assign img[ 8465] = 134;
assign img[ 8466] = 128;
assign img[ 8467] = 132;
assign img[ 8468] = 133;
assign img[ 8469] = 132;
assign img[ 8470] = 128;
assign img[ 8471] = 128;
assign img[ 8472] = 128;
assign img[ 8473] = 132;
assign img[ 8474] = 133;
assign img[ 8475] = 128;
assign img[ 8476] = 128;
assign img[ 8477] = 130;
assign img[ 8478] = 128;
assign img[ 8479] = 128;
assign img[ 8480] = 128;
assign img[ 8481] = 128;
assign img[ 8482] = 128;
assign img[ 8483] = 132;
assign img[ 8484] = 128;
assign img[ 8485] = 128;
assign img[ 8486] = 128;
assign img[ 8487] = 132;
assign img[ 8488] = 128;
assign img[ 8489] = 134;
assign img[ 8490] = 128;
assign img[ 8491] = 128;
assign img[ 8492] = 128;
assign img[ 8493] = 128;
assign img[ 8494] = 130;
assign img[ 8495] = 132;
assign img[ 8496] = 132;
assign img[ 8497] = 128;
assign img[ 8498] = 130;
assign img[ 8499] = 128;
assign img[ 8500] = 131;
assign img[ 8501] = 133;
assign img[ 8502] = 128;
assign img[ 8503] = 128;
assign img[ 8504] = 128;
assign img[ 8505] = 128;
assign img[ 8506] = 116;
assign img[ 8507] = 103;
assign img[ 8508] = 105;
assign img[ 8509] = 104;
assign img[ 8510] = 103;
assign img[ 8511] = 101;
assign img[ 8512] = 103;
assign img[ 8513] = 101;
assign img[ 8514] = 101;
assign img[ 8515] = 101;
assign img[ 8516] = 100;
assign img[ 8517] = 100;
assign img[ 8518] = 93;
assign img[ 8519] = 97;
assign img[ 8520] = 105;
assign img[ 8521] = 97;
assign img[ 8522] = 101;
assign img[ 8523] = 101;
assign img[ 8524] = 102;
assign img[ 8525] = 102;
assign img[ 8526] = 102;
assign img[ 8527] = 105;
assign img[ 8528] = 100;
assign img[ 8529] = 98;
assign img[ 8530] = 101;
assign img[ 8531] = 96;
assign img[ 8532] = 100;
assign img[ 8533] = 108;
assign img[ 8534] = 103;
assign img[ 8535] = 94;
assign img[ 8536] = 94;
assign img[ 8537] = 97;
assign img[ 8538] = 100;
assign img[ 8539] = 95;
assign img[ 8540] = 100;
assign img[ 8541] = 95;
assign img[ 8542] = 104;
assign img[ 8543] = 94;
assign img[ 8544] = 95;
assign img[ 8545] = 100;
assign img[ 8546] = 97;
assign img[ 8547] = 92;
assign img[ 8548] = 92;
assign img[ 8549] = 96;
assign img[ 8550] = 98;
assign img[ 8551] = 96;
assign img[ 8552] = 92;
assign img[ 8553] = 96;
assign img[ 8554] = 100;
assign img[ 8555] = 92;
assign img[ 8556] = 88;
assign img[ 8557] = 92;
assign img[ 8558] = 89;
assign img[ 8559] = 95;
assign img[ 8560] = 94;
assign img[ 8561] = 95;
assign img[ 8562] = 97;
assign img[ 8563] = 94;
assign img[ 8564] = 92;
assign img[ 8565] = 94;
assign img[ 8566] = 94;
assign img[ 8567] = 92;
assign img[ 8568] = 94;
assign img[ 8569] = 89;
assign img[ 8570] = 89;
assign img[ 8571] = 93;
assign img[ 8572] = 96;
assign img[ 8573] = 95;
assign img[ 8574] = 100;
assign img[ 8575] = 93;
assign img[ 8576] = 96;
assign img[ 8577] = 102;
assign img[ 8578] = 106;
assign img[ 8579] = 106;
assign img[ 8580] = 105;
assign img[ 8581] = 113;
assign img[ 8582] = 113;
assign img[ 8583] = 114;
assign img[ 8584] = 129;
assign img[ 8585] = 130;
assign img[ 8586] = 130;
assign img[ 8587] = 130;
assign img[ 8588] = 130;
assign img[ 8589] = 130;
assign img[ 8590] = 130;
assign img[ 8591] = 128;
assign img[ 8592] = 130;
assign img[ 8593] = 134;
assign img[ 8594] = 130;
assign img[ 8595] = 128;
assign img[ 8596] = 128;
assign img[ 8597] = 130;
assign img[ 8598] = 134;
assign img[ 8599] = 135;
assign img[ 8600] = 132;
assign img[ 8601] = 128;
assign img[ 8602] = 130;
assign img[ 8603] = 130;
assign img[ 8604] = 130;
assign img[ 8605] = 128;
assign img[ 8606] = 130;
assign img[ 8607] = 136;
assign img[ 8608] = 128;
assign img[ 8609] = 128;
assign img[ 8610] = 130;
assign img[ 8611] = 134;
assign img[ 8612] = 128;
assign img[ 8613] = 128;
assign img[ 8614] = 130;
assign img[ 8615] = 128;
assign img[ 8616] = 134;
assign img[ 8617] = 128;
assign img[ 8618] = 128;
assign img[ 8619] = 128;
assign img[ 8620] = 128;
assign img[ 8621] = 130;
assign img[ 8622] = 130;
assign img[ 8623] = 130;
assign img[ 8624] = 130;
assign img[ 8625] = 128;
assign img[ 8626] = 130;
assign img[ 8627] = 130;
assign img[ 8628] = 132;
assign img[ 8629] = 128;
assign img[ 8630] = 130;
assign img[ 8631] = 128;
assign img[ 8632] = 128;
assign img[ 8633] = 130;
assign img[ 8634] = 128;
assign img[ 8635] = 111;
assign img[ 8636] = 103;
assign img[ 8637] = 100;
assign img[ 8638] = 97;
assign img[ 8639] = 110;
assign img[ 8640] = 97;
assign img[ 8641] = 96;
assign img[ 8642] = 96;
assign img[ 8643] = 96;
assign img[ 8644] = 97;
assign img[ 8645] = 93;
assign img[ 8646] = 104;
assign img[ 8647] = 90;
assign img[ 8648] = 94;
assign img[ 8649] = 97;
assign img[ 8650] = 103;
assign img[ 8651] = 97;
assign img[ 8652] = 100;
assign img[ 8653] = 103;
assign img[ 8654] = 93;
assign img[ 8655] = 104;
assign img[ 8656] = 101;
assign img[ 8657] = 97;
assign img[ 8658] = 101;
assign img[ 8659] = 101;
assign img[ 8660] = 102;
assign img[ 8661] = 96;
assign img[ 8662] = 92;
assign img[ 8663] = 96;
assign img[ 8664] = 92;
assign img[ 8665] = 94;
assign img[ 8666] = 91;
assign img[ 8667] = 94;
assign img[ 8668] = 99;
assign img[ 8669] = 96;
assign img[ 8670] = 100;
assign img[ 8671] = 94;
assign img[ 8672] = 94;
assign img[ 8673] = 95;
assign img[ 8674] = 94;
assign img[ 8675] = 94;
assign img[ 8676] = 100;
assign img[ 8677] = 91;
assign img[ 8678] = 92;
assign img[ 8679] = 97;
assign img[ 8680] = 96;
assign img[ 8681] = 95;
assign img[ 8682] = 96;
assign img[ 8683] = 94;
assign img[ 8684] = 95;
assign img[ 8685] = 98;
assign img[ 8686] = 105;
assign img[ 8687] = 93;
assign img[ 8688] = 97;
assign img[ 8689] = 96;
assign img[ 8690] = 88;
assign img[ 8691] = 94;
assign img[ 8692] = 92;
assign img[ 8693] = 93;
assign img[ 8694] = 93;
assign img[ 8695] = 89;
assign img[ 8696] = 94;
assign img[ 8697] = 92;
assign img[ 8698] = 98;
assign img[ 8699] = 92;
assign img[ 8700] = 87;
assign img[ 8701] = 92;
assign img[ 8702] = 90;
assign img[ 8703] = 98;
assign img[ 8704] = 98;
assign img[ 8705] = 105;
assign img[ 8706] = 112;
assign img[ 8707] = 102;
assign img[ 8708] = 104;
assign img[ 8709] = 104;
assign img[ 8710] = 112;
assign img[ 8711] = 109;
assign img[ 8712] = 128;
assign img[ 8713] = 128;
assign img[ 8714] = 128;
assign img[ 8715] = 128;
assign img[ 8716] = 128;
assign img[ 8717] = 128;
assign img[ 8718] = 128;
assign img[ 8719] = 132;
assign img[ 8720] = 128;
assign img[ 8721] = 128;
assign img[ 8722] = 128;
assign img[ 8723] = 128;
assign img[ 8724] = 128;
assign img[ 8725] = 128;
assign img[ 8726] = 128;
assign img[ 8727] = 128;
assign img[ 8728] = 128;
assign img[ 8729] = 128;
assign img[ 8730] = 128;
assign img[ 8731] = 128;
assign img[ 8732] = 128;
assign img[ 8733] = 128;
assign img[ 8734] = 128;
assign img[ 8735] = 128;
assign img[ 8736] = 128;
assign img[ 8737] = 131;
assign img[ 8738] = 132;
assign img[ 8739] = 128;
assign img[ 8740] = 128;
assign img[ 8741] = 128;
assign img[ 8742] = 128;
assign img[ 8743] = 128;
assign img[ 8744] = 128;
assign img[ 8745] = 128;
assign img[ 8746] = 130;
assign img[ 8747] = 128;
assign img[ 8748] = 130;
assign img[ 8749] = 128;
assign img[ 8750] = 128;
assign img[ 8751] = 128;
assign img[ 8752] = 128;
assign img[ 8753] = 128;
assign img[ 8754] = 128;
assign img[ 8755] = 128;
assign img[ 8756] = 128;
assign img[ 8757] = 128;
assign img[ 8758] = 128;
assign img[ 8759] = 128;
assign img[ 8760] = 128;
assign img[ 8761] = 128;
assign img[ 8762] = 128;
assign img[ 8763] = 128;
assign img[ 8764] = 112;
assign img[ 8765] = 104;
assign img[ 8766] = 104;
assign img[ 8767] = 96;
assign img[ 8768] = 93;
assign img[ 8769] = 96;
assign img[ 8770] = 100;
assign img[ 8771] = 93;
assign img[ 8772] = 96;
assign img[ 8773] = 100;
assign img[ 8774] = 94;
assign img[ 8775] = 97;
assign img[ 8776] = 96;
assign img[ 8777] = 96;
assign img[ 8778] = 92;
assign img[ 8779] = 96;
assign img[ 8780] = 96;
assign img[ 8781] = 89;
assign img[ 8782] = 96;
assign img[ 8783] = 99;
assign img[ 8784] = 96;
assign img[ 8785] = 90;
assign img[ 8786] = 96;
assign img[ 8787] = 97;
assign img[ 8788] = 97;
assign img[ 8789] = 97;
assign img[ 8790] = 91;
assign img[ 8791] = 92;
assign img[ 8792] = 96;
assign img[ 8793] = 97;
assign img[ 8794] = 98;
assign img[ 8795] = 98;
assign img[ 8796] = 96;
assign img[ 8797] = 97;
assign img[ 8798] = 98;
assign img[ 8799] = 94;
assign img[ 8800] = 93;
assign img[ 8801] = 96;
assign img[ 8802] = 92;
assign img[ 8803] = 85;
assign img[ 8804] = 96;
assign img[ 8805] = 97;
assign img[ 8806] = 97;
assign img[ 8807] = 93;
assign img[ 8808] = 96;
assign img[ 8809] = 100;
assign img[ 8810] = 86;
assign img[ 8811] = 88;
assign img[ 8812] = 96;
assign img[ 8813] = 97;
assign img[ 8814] = 96;
assign img[ 8815] = 93;
assign img[ 8816] = 89;
assign img[ 8817] = 92;
assign img[ 8818] = 92;
assign img[ 8819] = 87;
assign img[ 8820] = 84;
assign img[ 8821] = 88;
assign img[ 8822] = 91;
assign img[ 8823] = 90;
assign img[ 8824] = 96;
assign img[ 8825] = 87;
assign img[ 8826] = 96;
assign img[ 8827] = 89;
assign img[ 8828] = 92;
assign img[ 8829] = 97;
assign img[ 8830] = 92;
assign img[ 8831] = 96;
assign img[ 8832] = 92;
assign img[ 8833] = 116;
assign img[ 8834] = 105;
assign img[ 8835] = 112;
assign img[ 8836] = 115;
assign img[ 8837] = 111;
assign img[ 8838] = 108;
assign img[ 8839] = 108;
assign img[ 8840] = 112;
assign img[ 8841] = 128;
assign img[ 8842] = 130;
assign img[ 8843] = 128;
assign img[ 8844] = 134;
assign img[ 8845] = 128;
assign img[ 8846] = 128;
assign img[ 8847] = 130;
assign img[ 8848] = 128;
assign img[ 8849] = 130;
assign img[ 8850] = 130;
assign img[ 8851] = 128;
assign img[ 8852] = 132;
assign img[ 8853] = 128;
assign img[ 8854] = 130;
assign img[ 8855] = 128;
assign img[ 8856] = 128;
assign img[ 8857] = 128;
assign img[ 8858] = 132;
assign img[ 8859] = 128;
assign img[ 8860] = 128;
assign img[ 8861] = 130;
assign img[ 8862] = 134;
assign img[ 8863] = 130;
assign img[ 8864] = 128;
assign img[ 8865] = 130;
assign img[ 8866] = 128;
assign img[ 8867] = 128;
assign img[ 8868] = 130;
assign img[ 8869] = 130;
assign img[ 8870] = 128;
assign img[ 8871] = 128;
assign img[ 8872] = 134;
assign img[ 8873] = 130;
assign img[ 8874] = 130;
assign img[ 8875] = 128;
assign img[ 8876] = 128;
assign img[ 8877] = 128;
assign img[ 8878] = 128;
assign img[ 8879] = 135;
assign img[ 8880] = 129;
assign img[ 8881] = 129;
assign img[ 8882] = 131;
assign img[ 8883] = 128;
assign img[ 8884] = 128;
assign img[ 8885] = 130;
assign img[ 8886] = 134;
assign img[ 8887] = 128;
assign img[ 8888] = 131;
assign img[ 8889] = 130;
assign img[ 8890] = 128;
assign img[ 8891] = 130;
assign img[ 8892] = 128;
assign img[ 8893] = 117;
assign img[ 8894] = 108;
assign img[ 8895] = 104;
assign img[ 8896] = 104;
assign img[ 8897] = 105;
assign img[ 8898] = 102;
assign img[ 8899] = 104;
assign img[ 8900] = 97;
assign img[ 8901] = 99;
assign img[ 8902] = 104;
assign img[ 8903] = 96;
assign img[ 8904] = 96;
assign img[ 8905] = 100;
assign img[ 8906] = 104;
assign img[ 8907] = 100;
assign img[ 8908] = 96;
assign img[ 8909] = 96;
assign img[ 8910] = 95;
assign img[ 8911] = 96;
assign img[ 8912] = 94;
assign img[ 8913] = 100;
assign img[ 8914] = 100;
assign img[ 8915] = 104;
assign img[ 8916] = 100;
assign img[ 8917] = 104;
assign img[ 8918] = 96;
assign img[ 8919] = 98;
assign img[ 8920] = 96;
assign img[ 8921] = 100;
assign img[ 8922] = 97;
assign img[ 8923] = 98;
assign img[ 8924] = 97;
assign img[ 8925] = 100;
assign img[ 8926] = 100;
assign img[ 8927] = 97;
assign img[ 8928] = 92;
assign img[ 8929] = 96;
assign img[ 8930] = 97;
assign img[ 8931] = 95;
assign img[ 8932] = 92;
assign img[ 8933] = 96;
assign img[ 8934] = 102;
assign img[ 8935] = 98;
assign img[ 8936] = 94;
assign img[ 8937] = 96;
assign img[ 8938] = 104;
assign img[ 8939] = 93;
assign img[ 8940] = 95;
assign img[ 8941] = 100;
assign img[ 8942] = 92;
assign img[ 8943] = 92;
assign img[ 8944] = 96;
assign img[ 8945] = 97;
assign img[ 8946] = 96;
assign img[ 8947] = 94;
assign img[ 8948] = 100;
assign img[ 8949] = 93;
assign img[ 8950] = 97;
assign img[ 8951] = 102;
assign img[ 8952] = 96;
assign img[ 8953] = 94;
assign img[ 8954] = 94;
assign img[ 8955] = 93;
assign img[ 8956] = 92;
assign img[ 8957] = 97;
assign img[ 8958] = 85;
assign img[ 8959] = 94;
assign img[ 8960] = 98;
assign img[ 8961] = 83;
assign img[ 8962] = 84;
assign img[ 8963] = 76;
assign img[ 8964] = 72;
assign img[ 8965] = 83;
assign img[ 8966] = 73;
assign img[ 8967] = 78;
assign img[ 8968] = 92;
assign img[ 8969] = 88;
assign img[ 8970] = 99;
assign img[ 8971] = 96;
assign img[ 8972] = 108;
assign img[ 8973] = 99;
assign img[ 8974] = 94;
assign img[ 8975] = 100;
assign img[ 8976] = 100;
assign img[ 8977] = 102;
assign img[ 8978] = 102;
assign img[ 8979] = 104;
assign img[ 8980] = 104;
assign img[ 8981] = 100;
assign img[ 8982] = 100;
assign img[ 8983] = 96;
assign img[ 8984] = 100;
assign img[ 8985] = 104;
assign img[ 8986] = 102;
assign img[ 8987] = 98;
assign img[ 8988] = 103;
assign img[ 8989] = 99;
assign img[ 8990] = 96;
assign img[ 8991] = 102;
assign img[ 8992] = 106;
assign img[ 8993] = 99;
assign img[ 8994] = 103;
assign img[ 8995] = 100;
assign img[ 8996] = 102;
assign img[ 8997] = 96;
assign img[ 8998] = 100;
assign img[ 8999] = 99;
assign img[ 9000] = 97;
assign img[ 9001] = 98;
assign img[ 9002] = 102;
assign img[ 9003] = 104;
assign img[ 9004] = 104;
assign img[ 9005] = 100;
assign img[ 9006] = 97;
assign img[ 9007] = 98;
assign img[ 9008] = 101;
assign img[ 9009] = 98;
assign img[ 9010] = 98;
assign img[ 9011] = 97;
assign img[ 9012] = 106;
assign img[ 9013] = 98;
assign img[ 9014] = 98;
assign img[ 9015] = 97;
assign img[ 9016] = 105;
assign img[ 9017] = 100;
assign img[ 9018] = 100;
assign img[ 9019] = 108;
assign img[ 9020] = 99;
assign img[ 9021] = 89;
assign img[ 9022] = 96;
assign img[ 9023] = 89;
assign img[ 9024] = 85;
assign img[ 9025] = 75;
assign img[ 9026] = 79;
assign img[ 9027] = 83;
assign img[ 9028] = 72;
assign img[ 9029] = 83;
assign img[ 9030] = 73;
assign img[ 9031] = 78;
assign img[ 9032] = 73;
assign img[ 9033] = 74;
assign img[ 9034] = 71;
assign img[ 9035] = 73;
assign img[ 9036] = 76;
assign img[ 9037] = 69;
assign img[ 9038] = 77;
assign img[ 9039] = 68;
assign img[ 9040] = 68;
assign img[ 9041] = 68;
assign img[ 9042] = 68;
assign img[ 9043] = 69;
assign img[ 9044] = 70;
assign img[ 9045] = 70;
assign img[ 9046] = 65;
assign img[ 9047] = 70;
assign img[ 9048] = 70;
assign img[ 9049] = 72;
assign img[ 9050] = 71;
assign img[ 9051] = 74;
assign img[ 9052] = 71;
assign img[ 9053] = 65;
assign img[ 9054] = 71;
assign img[ 9055] = 73;
assign img[ 9056] = 69;
assign img[ 9057] = 70;
assign img[ 9058] = 72;
assign img[ 9059] = 70;
assign img[ 9060] = 69;
assign img[ 9061] = 72;
assign img[ 9062] = 73;
assign img[ 9063] = 72;
assign img[ 9064] = 73;
assign img[ 9065] = 72;
assign img[ 9066] = 68;
assign img[ 9067] = 64;
assign img[ 9068] = 66;
assign img[ 9069] = 66;
assign img[ 9070] = 69;
assign img[ 9071] = 69;
assign img[ 9072] = 71;
assign img[ 9073] = 66;
assign img[ 9074] = 71;
assign img[ 9075] = 70;
assign img[ 9076] = 64;
assign img[ 9077] = 70;
assign img[ 9078] = 73;
assign img[ 9079] = 70;
assign img[ 9080] = 66;
assign img[ 9081] = 71;
assign img[ 9082] = 73;
assign img[ 9083] = 68;
assign img[ 9084] = 72;
assign img[ 9085] = 73;
assign img[ 9086] = 71;
assign img[ 9087] = 70;
assign img[ 9088] = 64;
assign img[ 9089] = 97;
assign img[ 9090] = 96;
assign img[ 9091] = 94;
assign img[ 9092] = 92;
assign img[ 9093] = 94;
assign img[ 9094] = 93;
assign img[ 9095] = 97;
assign img[ 9096] = 96;
assign img[ 9097] = 105;
assign img[ 9098] = 128;
assign img[ 9099] = 110;
assign img[ 9100] = 109;
assign img[ 9101] = 105;
assign img[ 9102] = 113;
assign img[ 9103] = 113;
assign img[ 9104] = 113;
assign img[ 9105] = 109;
assign img[ 9106] = 128;
assign img[ 9107] = 117;
assign img[ 9108] = 112;
assign img[ 9109] = 108;
assign img[ 9110] = 107;
assign img[ 9111] = 120;
assign img[ 9112] = 117;
assign img[ 9113] = 113;
assign img[ 9114] = 117;
assign img[ 9115] = 109;
assign img[ 9116] = 110;
assign img[ 9117] = 113;
assign img[ 9118] = 105;
assign img[ 9119] = 108;
assign img[ 9120] = 104;
assign img[ 9121] = 117;
assign img[ 9122] = 109;
assign img[ 9123] = 114;
assign img[ 9124] = 106;
assign img[ 9125] = 110;
assign img[ 9126] = 117;
assign img[ 9127] = 105;
assign img[ 9128] = 104;
assign img[ 9129] = 113;
assign img[ 9130] = 110;
assign img[ 9131] = 113;
assign img[ 9132] = 113;
assign img[ 9133] = 110;
assign img[ 9134] = 117;
assign img[ 9135] = 113;
assign img[ 9136] = 109;
assign img[ 9137] = 105;
assign img[ 9138] = 117;
assign img[ 9139] = 117;
assign img[ 9140] = 108;
assign img[ 9141] = 113;
assign img[ 9142] = 112;
assign img[ 9143] = 105;
assign img[ 9144] = 113;
assign img[ 9145] = 117;
assign img[ 9146] = 111;
assign img[ 9147] = 113;
assign img[ 9148] = 109;
assign img[ 9149] = 109;
assign img[ 9150] = 101;
assign img[ 9151] = 105;
assign img[ 9152] = 97;
assign img[ 9153] = 96;
assign img[ 9154] = 94;
assign img[ 9155] = 96;
assign img[ 9156] = 85;
assign img[ 9157] = 89;
assign img[ 9158] = 89;
assign img[ 9159] = 93;
assign img[ 9160] = 85;
assign img[ 9161] = 86;
assign img[ 9162] = 88;
assign img[ 9163] = 89;
assign img[ 9164] = 89;
assign img[ 9165] = 89;
assign img[ 9166] = 85;
assign img[ 9167] = 85;
assign img[ 9168] = 77;
assign img[ 9169] = 82;
assign img[ 9170] = 82;
assign img[ 9171] = 88;
assign img[ 9172] = 87;
assign img[ 9173] = 80;
assign img[ 9174] = 90;
assign img[ 9175] = 92;
assign img[ 9176] = 84;
assign img[ 9177] = 85;
assign img[ 9178] = 84;
assign img[ 9179] = 84;
assign img[ 9180] = 80;
assign img[ 9181] = 77;
assign img[ 9182] = 80;
assign img[ 9183] = 77;
assign img[ 9184] = 84;
assign img[ 9185] = 92;
assign img[ 9186] = 77;
assign img[ 9187] = 85;
assign img[ 9188] = 84;
assign img[ 9189] = 85;
assign img[ 9190] = 79;
assign img[ 9191] = 81;
assign img[ 9192] = 84;
assign img[ 9193] = 78;
assign img[ 9194] = 89;
assign img[ 9195] = 87;
assign img[ 9196] = 76;
assign img[ 9197] = 77;
assign img[ 9198] = 85;
assign img[ 9199] = 76;
assign img[ 9200] = 78;
assign img[ 9201] = 77;
assign img[ 9202] = 79;
assign img[ 9203] = 80;
assign img[ 9204] = 79;
assign img[ 9205] = 81;
assign img[ 9206] = 79;
assign img[ 9207] = 72;
assign img[ 9208] = 84;
assign img[ 9209] = 85;
assign img[ 9210] = 76;
assign img[ 9211] = 74;
assign img[ 9212] = 86;
assign img[ 9213] = 84;
assign img[ 9214] = 77;
assign img[ 9215] = 81;
assign img[ 9216] = 79;
assign img[ 9217] = 84;
assign img[ 9218] = 77;
assign img[ 9219] = 80;
assign img[ 9220] = 80;
assign img[ 9221] = 80;
assign img[ 9222] = 85;
assign img[ 9223] = 81;
assign img[ 9224] = 88;
assign img[ 9225] = 94;
assign img[ 9226] = 100;
assign img[ 9227] = 100;
assign img[ 9228] = 98;
assign img[ 9229] = 98;
assign img[ 9230] = 105;
assign img[ 9231] = 105;
assign img[ 9232] = 101;
assign img[ 9233] = 97;
assign img[ 9234] = 102;
assign img[ 9235] = 101;
assign img[ 9236] = 101;
assign img[ 9237] = 100;
assign img[ 9238] = 97;
assign img[ 9239] = 101;
assign img[ 9240] = 104;
assign img[ 9241] = 102;
assign img[ 9242] = 106;
assign img[ 9243] = 108;
assign img[ 9244] = 97;
assign img[ 9245] = 101;
assign img[ 9246] = 98;
assign img[ 9247] = 104;
assign img[ 9248] = 111;
assign img[ 9249] = 97;
assign img[ 9250] = 96;
assign img[ 9251] = 102;
assign img[ 9252] = 107;
assign img[ 9253] = 101;
assign img[ 9254] = 96;
assign img[ 9255] = 113;
assign img[ 9256] = 102;
assign img[ 9257] = 97;
assign img[ 9258] = 105;
assign img[ 9259] = 100;
assign img[ 9260] = 97;
assign img[ 9261] = 100;
assign img[ 9262] = 100;
assign img[ 9263] = 104;
assign img[ 9264] = 101;
assign img[ 9265] = 103;
assign img[ 9266] = 103;
assign img[ 9267] = 101;
assign img[ 9268] = 96;
assign img[ 9269] = 96;
assign img[ 9270] = 97;
assign img[ 9271] = 104;
assign img[ 9272] = 110;
assign img[ 9273] = 105;
assign img[ 9274] = 96;
assign img[ 9275] = 96;
assign img[ 9276] = 105;
assign img[ 9277] = 97;
assign img[ 9278] = 98;
assign img[ 9279] = 96;
assign img[ 9280] = 92;
assign img[ 9281] = 89;
assign img[ 9282] = 77;
assign img[ 9283] = 86;
assign img[ 9284] = 77;
assign img[ 9285] = 78;
assign img[ 9286] = 80;
assign img[ 9287] = 75;
assign img[ 9288] = 76;
assign img[ 9289] = 84;
assign img[ 9290] = 73;
assign img[ 9291] = 69;
assign img[ 9292] = 64;
assign img[ 9293] = 76;
assign img[ 9294] = 74;
assign img[ 9295] = 78;
assign img[ 9296] = 78;
assign img[ 9297] = 71;
assign img[ 9298] = 68;
assign img[ 9299] = 69;
assign img[ 9300] = 73;
assign img[ 9301] = 68;
assign img[ 9302] = 73;
assign img[ 9303] = 76;
assign img[ 9304] = 76;
assign img[ 9305] = 68;
assign img[ 9306] = 77;
assign img[ 9307] = 71;
assign img[ 9308] = 72;
assign img[ 9309] = 72;
assign img[ 9310] = 80;
assign img[ 9311] = 70;
assign img[ 9312] = 71;
assign img[ 9313] = 70;
assign img[ 9314] = 71;
assign img[ 9315] = 77;
assign img[ 9316] = 76;
assign img[ 9317] = 72;
assign img[ 9318] = 77;
assign img[ 9319] = 73;
assign img[ 9320] = 69;
assign img[ 9321] = 71;
assign img[ 9322] = 76;
assign img[ 9323] = 71;
assign img[ 9324] = 71;
assign img[ 9325] = 74;
assign img[ 9326] = 76;
assign img[ 9327] = 68;
assign img[ 9328] = 68;
assign img[ 9329] = 66;
assign img[ 9330] = 70;
assign img[ 9331] = 78;
assign img[ 9332] = 68;
assign img[ 9333] = 73;
assign img[ 9334] = 76;
assign img[ 9335] = 65;
assign img[ 9336] = 72;
assign img[ 9337] = 76;
assign img[ 9338] = 66;
assign img[ 9339] = 70;
assign img[ 9340] = 69;
assign img[ 9341] = 68;
assign img[ 9342] = 71;
assign img[ 9343] = 71;
assign img[ 9344] = 72;
assign img[ 9345] = 79;
assign img[ 9346] = 74;
assign img[ 9347] = 81;
assign img[ 9348] = 76;
assign img[ 9349] = 76;
assign img[ 9350] = 80;
assign img[ 9351] = 76;
assign img[ 9352] = 85;
assign img[ 9353] = 92;
assign img[ 9354] = 91;
assign img[ 9355] = 101;
assign img[ 9356] = 96;
assign img[ 9357] = 93;
assign img[ 9358] = 94;
assign img[ 9359] = 94;
assign img[ 9360] = 94;
assign img[ 9361] = 95;
assign img[ 9362] = 93;
assign img[ 9363] = 97;
assign img[ 9364] = 90;
assign img[ 9365] = 96;
assign img[ 9366] = 95;
assign img[ 9367] = 92;
assign img[ 9368] = 94;
assign img[ 9369] = 89;
assign img[ 9370] = 94;
assign img[ 9371] = 86;
assign img[ 9372] = 96;
assign img[ 9373] = 96;
assign img[ 9374] = 95;
assign img[ 9375] = 96;
assign img[ 9376] = 93;
assign img[ 9377] = 97;
assign img[ 9378] = 95;
assign img[ 9379] = 92;
assign img[ 9380] = 95;
assign img[ 9381] = 93;
assign img[ 9382] = 94;
assign img[ 9383] = 88;
assign img[ 9384] = 92;
assign img[ 9385] = 93;
assign img[ 9386] = 92;
assign img[ 9387] = 91;
assign img[ 9388] = 94;
assign img[ 9389] = 84;
assign img[ 9390] = 102;
assign img[ 9391] = 96;
assign img[ 9392] = 92;
assign img[ 9393] = 96;
assign img[ 9394] = 89;
assign img[ 9395] = 100;
assign img[ 9396] = 94;
assign img[ 9397] = 92;
assign img[ 9398] = 100;
assign img[ 9399] = 91;
assign img[ 9400] = 93;
assign img[ 9401] = 92;
assign img[ 9402] = 88;
assign img[ 9403] = 96;
assign img[ 9404] = 88;
assign img[ 9405] = 86;
assign img[ 9406] = 89;
assign img[ 9407] = 92;
assign img[ 9408] = 87;
assign img[ 9409] = 86;
assign img[ 9410] = 78;
assign img[ 9411] = 78;
assign img[ 9412] = 69;
assign img[ 9413] = 72;
assign img[ 9414] = 72;
assign img[ 9415] = 69;
assign img[ 9416] = 68;
assign img[ 9417] = 73;
assign img[ 9418] = 76;
assign img[ 9419] = 70;
assign img[ 9420] = 65;
assign img[ 9421] = 64;
assign img[ 9422] = 70;
assign img[ 9423] = 71;
assign img[ 9424] = 68;
assign img[ 9425] = 58;
assign img[ 9426] = 65;
assign img[ 9427] = 64;
assign img[ 9428] = 65;
assign img[ 9429] = 65;
assign img[ 9430] = 68;
assign img[ 9431] = 70;
assign img[ 9432] = 64;
assign img[ 9433] = 64;
assign img[ 9434] = 68;
assign img[ 9435] = 68;
assign img[ 9436] = 64;
assign img[ 9437] = 68;
assign img[ 9438] = 70;
assign img[ 9439] = 70;
assign img[ 9440] = 64;
assign img[ 9441] = 66;
assign img[ 9442] = 64;
assign img[ 9443] = 64;
assign img[ 9444] = 64;
assign img[ 9445] = 70;
assign img[ 9446] = 64;
assign img[ 9447] = 68;
assign img[ 9448] = 68;
assign img[ 9449] = 72;
assign img[ 9450] = 68;
assign img[ 9451] = 70;
assign img[ 9452] = 69;
assign img[ 9453] = 64;
assign img[ 9454] = 64;
assign img[ 9455] = 70;
assign img[ 9456] = 64;
assign img[ 9457] = 66;
assign img[ 9458] = 68;
assign img[ 9459] = 64;
assign img[ 9460] = 64;
assign img[ 9461] = 64;
assign img[ 9462] = 66;
assign img[ 9463] = 64;
assign img[ 9464] = 64;
assign img[ 9465] = 64;
assign img[ 9466] = 70;
assign img[ 9467] = 64;
assign img[ 9468] = 64;
assign img[ 9469] = 60;
assign img[ 9470] = 65;
assign img[ 9471] = 66;
assign img[ 9472] = 64;
assign img[ 9473] = 96;
assign img[ 9474] = 94;
assign img[ 9475] = 92;
assign img[ 9476] = 83;
assign img[ 9477] = 86;
assign img[ 9478] = 99;
assign img[ 9479] = 100;
assign img[ 9480] = 100;
assign img[ 9481] = 106;
assign img[ 9482] = 109;
assign img[ 9483] = 101;
assign img[ 9484] = 108;
assign img[ 9485] = 128;
assign img[ 9486] = 96;
assign img[ 9487] = 107;
assign img[ 9488] = 109;
assign img[ 9489] = 106;
assign img[ 9490] = 110;
assign img[ 9491] = 104;
assign img[ 9492] = 101;
assign img[ 9493] = 108;
assign img[ 9494] = 103;
assign img[ 9495] = 104;
assign img[ 9496] = 108;
assign img[ 9497] = 104;
assign img[ 9498] = 105;
assign img[ 9499] = 111;
assign img[ 9500] = 104;
assign img[ 9501] = 109;
assign img[ 9502] = 109;
assign img[ 9503] = 104;
assign img[ 9504] = 113;
assign img[ 9505] = 105;
assign img[ 9506] = 104;
assign img[ 9507] = 108;
assign img[ 9508] = 105;
assign img[ 9509] = 97;
assign img[ 9510] = 110;
assign img[ 9511] = 100;
assign img[ 9512] = 104;
assign img[ 9513] = 106;
assign img[ 9514] = 104;
assign img[ 9515] = 108;
assign img[ 9516] = 101;
assign img[ 9517] = 102;
assign img[ 9518] = 106;
assign img[ 9519] = 107;
assign img[ 9520] = 108;
assign img[ 9521] = 104;
assign img[ 9522] = 109;
assign img[ 9523] = 100;
assign img[ 9524] = 100;
assign img[ 9525] = 106;
assign img[ 9526] = 101;
assign img[ 9527] = 102;
assign img[ 9528] = 104;
assign img[ 9529] = 108;
assign img[ 9530] = 106;
assign img[ 9531] = 102;
assign img[ 9532] = 105;
assign img[ 9533] = 99;
assign img[ 9534] = 106;
assign img[ 9535] = 101;
assign img[ 9536] = 97;
assign img[ 9537] = 100;
assign img[ 9538] = 96;
assign img[ 9539] = 90;
assign img[ 9540] = 81;
assign img[ 9541] = 84;
assign img[ 9542] = 89;
assign img[ 9543] = 78;
assign img[ 9544] = 82;
assign img[ 9545] = 87;
assign img[ 9546] = 80;
assign img[ 9547] = 81;
assign img[ 9548] = 82;
assign img[ 9549] = 84;
assign img[ 9550] = 73;
assign img[ 9551] = 81;
assign img[ 9552] = 81;
assign img[ 9553] = 80;
assign img[ 9554] = 73;
assign img[ 9555] = 82;
assign img[ 9556] = 80;
assign img[ 9557] = 72;
assign img[ 9558] = 73;
assign img[ 9559] = 80;
assign img[ 9560] = 81;
assign img[ 9561] = 69;
assign img[ 9562] = 72;
assign img[ 9563] = 80;
assign img[ 9564] = 86;
assign img[ 9565] = 76;
assign img[ 9566] = 81;
assign img[ 9567] = 73;
assign img[ 9568] = 81;
assign img[ 9569] = 82;
assign img[ 9570] = 80;
assign img[ 9571] = 73;
assign img[ 9572] = 79;
assign img[ 9573] = 81;
assign img[ 9574] = 77;
assign img[ 9575] = 82;
assign img[ 9576] = 81;
assign img[ 9577] = 73;
assign img[ 9578] = 81;
assign img[ 9579] = 82;
assign img[ 9580] = 82;
assign img[ 9581] = 76;
assign img[ 9582] = 81;
assign img[ 9583] = 81;
assign img[ 9584] = 73;
assign img[ 9585] = 82;
assign img[ 9586] = 77;
assign img[ 9587] = 72;
assign img[ 9588] = 84;
assign img[ 9589] = 74;
assign img[ 9590] = 72;
assign img[ 9591] = 70;
assign img[ 9592] = 77;
assign img[ 9593] = 82;
assign img[ 9594] = 76;
assign img[ 9595] = 81;
assign img[ 9596] = 66;
assign img[ 9597] = 70;
assign img[ 9598] = 73;
assign img[ 9599] = 73;
assign img[ 9600] = 80;
assign img[ 9601] = 54;
assign img[ 9602] = 64;
assign img[ 9603] = 58;
assign img[ 9604] = 64;
assign img[ 9605] = 64;
assign img[ 9606] = 56;
assign img[ 9607] = 67;
assign img[ 9608] = 72;
assign img[ 9609] = 73;
assign img[ 9610] = 80;
assign img[ 9611] = 73;
assign img[ 9612] = 69;
assign img[ 9613] = 76;
assign img[ 9614] = 80;
assign img[ 9615] = 66;
assign img[ 9616] = 74;
assign img[ 9617] = 73;
assign img[ 9618] = 72;
assign img[ 9619] = 69;
assign img[ 9620] = 73;
assign img[ 9621] = 69;
assign img[ 9622] = 72;
assign img[ 9623] = 81;
assign img[ 9624] = 73;
assign img[ 9625] = 76;
assign img[ 9626] = 70;
assign img[ 9627] = 77;
assign img[ 9628] = 77;
assign img[ 9629] = 74;
assign img[ 9630] = 69;
assign img[ 9631] = 83;
assign img[ 9632] = 73;
assign img[ 9633] = 73;
assign img[ 9634] = 73;
assign img[ 9635] = 73;
assign img[ 9636] = 77;
assign img[ 9637] = 74;
assign img[ 9638] = 81;
assign img[ 9639] = 77;
assign img[ 9640] = 80;
assign img[ 9641] = 73;
assign img[ 9642] = 73;
assign img[ 9643] = 80;
assign img[ 9644] = 66;
assign img[ 9645] = 72;
assign img[ 9646] = 67;
assign img[ 9647] = 82;
assign img[ 9648] = 74;
assign img[ 9649] = 76;
assign img[ 9650] = 78;
assign img[ 9651] = 75;
assign img[ 9652] = 77;
assign img[ 9653] = 69;
assign img[ 9654] = 76;
assign img[ 9655] = 74;
assign img[ 9656] = 80;
assign img[ 9657] = 74;
assign img[ 9658] = 72;
assign img[ 9659] = 74;
assign img[ 9660] = 73;
assign img[ 9661] = 73;
assign img[ 9662] = 76;
assign img[ 9663] = 80;
assign img[ 9664] = 74;
assign img[ 9665] = 75;
assign img[ 9666] = 65;
assign img[ 9667] = 66;
assign img[ 9668] = 64;
assign img[ 9669] = 53;
assign img[ 9670] = 54;
assign img[ 9671] = 51;
assign img[ 9672] = 56;
assign img[ 9673] = 56;
assign img[ 9674] = 53;
assign img[ 9675] = 50;
assign img[ 9676] = 54;
assign img[ 9677] = 53;
assign img[ 9678] = 50;
assign img[ 9679] = 50;
assign img[ 9680] = 48;
assign img[ 9681] = 50;
assign img[ 9682] = 54;
assign img[ 9683] = 54;
assign img[ 9684] = 54;
assign img[ 9685] = 49;
assign img[ 9686] = 49;
assign img[ 9687] = 48;
assign img[ 9688] = 46;
assign img[ 9689] = 48;
assign img[ 9690] = 48;
assign img[ 9691] = 46;
assign img[ 9692] = 49;
assign img[ 9693] = 52;
assign img[ 9694] = 46;
assign img[ 9695] = 44;
assign img[ 9696] = 53;
assign img[ 9697] = 48;
assign img[ 9698] = 55;
assign img[ 9699] = 53;
assign img[ 9700] = 42;
assign img[ 9701] = 55;
assign img[ 9702] = 54;
assign img[ 9703] = 45;
assign img[ 9704] = 50;
assign img[ 9705] = 48;
assign img[ 9706] = 49;
assign img[ 9707] = 54;
assign img[ 9708] = 46;
assign img[ 9709] = 49;
assign img[ 9710] = 46;
assign img[ 9711] = 46;
assign img[ 9712] = 43;
assign img[ 9713] = 51;
assign img[ 9714] = 55;
assign img[ 9715] = 47;
assign img[ 9716] = 44;
assign img[ 9717] = 39;
assign img[ 9718] = 47;
assign img[ 9719] = 46;
assign img[ 9720] = 49;
assign img[ 9721] = 42;
assign img[ 9722] = 48;
assign img[ 9723] = 49;
assign img[ 9724] = 44;
assign img[ 9725] = 47;
assign img[ 9726] = 44;
assign img[ 9727] = 58;
assign img[ 9728] = 47;
assign img[ 9729] = 69;
assign img[ 9730] = 62;
assign img[ 9731] = 64;
assign img[ 9732] = 66;
assign img[ 9733] = 64;
assign img[ 9734] = 72;
assign img[ 9735] = 74;
assign img[ 9736] = 74;
assign img[ 9737] = 80;
assign img[ 9738] = 85;
assign img[ 9739] = 81;
assign img[ 9740] = 90;
assign img[ 9741] = 81;
assign img[ 9742] = 89;
assign img[ 9743] = 81;
assign img[ 9744] = 85;
assign img[ 9745] = 82;
assign img[ 9746] = 80;
assign img[ 9747] = 88;
assign img[ 9748] = 93;
assign img[ 9749] = 81;
assign img[ 9750] = 84;
assign img[ 9751] = 96;
assign img[ 9752] = 84;
assign img[ 9753] = 86;
assign img[ 9754] = 89;
assign img[ 9755] = 89;
assign img[ 9756] = 81;
assign img[ 9757] = 82;
assign img[ 9758] = 88;
assign img[ 9759] = 89;
assign img[ 9760] = 88;
assign img[ 9761] = 89;
assign img[ 9762] = 82;
assign img[ 9763] = 92;
assign img[ 9764] = 81;
assign img[ 9765] = 82;
assign img[ 9766] = 81;
assign img[ 9767] = 77;
assign img[ 9768] = 85;
assign img[ 9769] = 84;
assign img[ 9770] = 85;
assign img[ 9771] = 96;
assign img[ 9772] = 94;
assign img[ 9773] = 89;
assign img[ 9774] = 84;
assign img[ 9775] = 86;
assign img[ 9776] = 90;
assign img[ 9777] = 88;
assign img[ 9778] = 88;
assign img[ 9779] = 87;
assign img[ 9780] = 81;
assign img[ 9781] = 85;
assign img[ 9782] = 96;
assign img[ 9783] = 84;
assign img[ 9784] = 86;
assign img[ 9785] = 84;
assign img[ 9786] = 85;
assign img[ 9787] = 92;
assign img[ 9788] = 97;
assign img[ 9789] = 86;
assign img[ 9790] = 84;
assign img[ 9791] = 87;
assign img[ 9792] = 89;
assign img[ 9793] = 85;
assign img[ 9794] = 86;
assign img[ 9795] = 77;
assign img[ 9796] = 69;
assign img[ 9797] = 67;
assign img[ 9798] = 66;
assign img[ 9799] = 64;
assign img[ 9800] = 65;
assign img[ 9801] = 64;
assign img[ 9802] = 64;
assign img[ 9803] = 58;
assign img[ 9804] = 68;
assign img[ 9805] = 58;
assign img[ 9806] = 64;
assign img[ 9807] = 70;
assign img[ 9808] = 60;
assign img[ 9809] = 56;
assign img[ 9810] = 64;
assign img[ 9811] = 64;
assign img[ 9812] = 64;
assign img[ 9813] = 59;
assign img[ 9814] = 64;
assign img[ 9815] = 60;
assign img[ 9816] = 54;
assign img[ 9817] = 64;
assign img[ 9818] = 64;
assign img[ 9819] = 64;
assign img[ 9820] = 56;
assign img[ 9821] = 64;
assign img[ 9822] = 56;
assign img[ 9823] = 64;
assign img[ 9824] = 64;
assign img[ 9825] = 58;
assign img[ 9826] = 56;
assign img[ 9827] = 64;
assign img[ 9828] = 54;
assign img[ 9829] = 64;
assign img[ 9830] = 59;
assign img[ 9831] = 56;
assign img[ 9832] = 55;
assign img[ 9833] = 46;
assign img[ 9834] = 64;
assign img[ 9835] = 56;
assign img[ 9836] = 64;
assign img[ 9837] = 64;
assign img[ 9838] = 64;
assign img[ 9839] = 64;
assign img[ 9840] = 56;
assign img[ 9841] = 64;
assign img[ 9842] = 64;
assign img[ 9843] = 64;
assign img[ 9844] = 55;
assign img[ 9845] = 64;
assign img[ 9846] = 54;
assign img[ 9847] = 56;
assign img[ 9848] = 53;
assign img[ 9849] = 55;
assign img[ 9850] = 64;
assign img[ 9851] = 53;
assign img[ 9852] = 55;
assign img[ 9853] = 64;
assign img[ 9854] = 56;
assign img[ 9855] = 55;
assign img[ 9856] = 60;
assign img[ 9857] = 69;
assign img[ 9858] = 68;
assign img[ 9859] = 78;
assign img[ 9860] = 64;
assign img[ 9861] = 71;
assign img[ 9862] = 72;
assign img[ 9863] = 72;
assign img[ 9864] = 80;
assign img[ 9865] = 85;
assign img[ 9866] = 92;
assign img[ 9867] = 87;
assign img[ 9868] = 90;
assign img[ 9869] = 85;
assign img[ 9870] = 85;
assign img[ 9871] = 91;
assign img[ 9872] = 80;
assign img[ 9873] = 89;
assign img[ 9874] = 88;
assign img[ 9875] = 89;
assign img[ 9876] = 89;
assign img[ 9877] = 90;
assign img[ 9878] = 97;
assign img[ 9879] = 86;
assign img[ 9880] = 88;
assign img[ 9881] = 96;
assign img[ 9882] = 93;
assign img[ 9883] = 97;
assign img[ 9884] = 90;
assign img[ 9885] = 92;
assign img[ 9886] = 93;
assign img[ 9887] = 96;
assign img[ 9888] = 85;
assign img[ 9889] = 89;
assign img[ 9890] = 97;
assign img[ 9891] = 97;
assign img[ 9892] = 93;
assign img[ 9893] = 96;
assign img[ 9894] = 89;
assign img[ 9895] = 97;
assign img[ 9896] = 90;
assign img[ 9897] = 89;
assign img[ 9898] = 97;
assign img[ 9899] = 91;
assign img[ 9900] = 96;
assign img[ 9901] = 96;
assign img[ 9902] = 89;
assign img[ 9903] = 97;
assign img[ 9904] = 96;
assign img[ 9905] = 92;
assign img[ 9906] = 89;
assign img[ 9907] = 96;
assign img[ 9908] = 88;
assign img[ 9909] = 93;
assign img[ 9910] = 89;
assign img[ 9911] = 90;
assign img[ 9912] = 89;
assign img[ 9913] = 97;
assign img[ 9914] = 89;
assign img[ 9915] = 90;
assign img[ 9916] = 90;
assign img[ 9917] = 92;
assign img[ 9918] = 89;
assign img[ 9919] = 85;
assign img[ 9920] = 82;
assign img[ 9921] = 89;
assign img[ 9922] = 82;
assign img[ 9923] = 85;
assign img[ 9924] = 81;
assign img[ 9925] = 81;
assign img[ 9926] = 72;
assign img[ 9927] = 65;
assign img[ 9928] = 64;
assign img[ 9929] = 73;
assign img[ 9930] = 60;
assign img[ 9931] = 65;
assign img[ 9932] = 65;
assign img[ 9933] = 64;
assign img[ 9934] = 66;
assign img[ 9935] = 66;
assign img[ 9936] = 58;
assign img[ 9937] = 64;
assign img[ 9938] = 64;
assign img[ 9939] = 66;
assign img[ 9940] = 64;
assign img[ 9941] = 64;
assign img[ 9942] = 64;
assign img[ 9943] = 56;
assign img[ 9944] = 64;
assign img[ 9945] = 64;
assign img[ 9946] = 64;
assign img[ 9947] = 64;
assign img[ 9948] = 50;
assign img[ 9949] = 64;
assign img[ 9950] = 64;
assign img[ 9951] = 60;
assign img[ 9952] = 64;
assign img[ 9953] = 59;
assign img[ 9954] = 64;
assign img[ 9955] = 64;
assign img[ 9956] = 64;
assign img[ 9957] = 64;
assign img[ 9958] = 66;
assign img[ 9959] = 57;
assign img[ 9960] = 58;
assign img[ 9961] = 64;
assign img[ 9962] = 60;
assign img[ 9963] = 64;
assign img[ 9964] = 56;
assign img[ 9965] = 56;
assign img[ 9966] = 64;
assign img[ 9967] = 65;
assign img[ 9968] = 64;
assign img[ 9969] = 66;
assign img[ 9970] = 64;
assign img[ 9971] = 59;
assign img[ 9972] = 64;
assign img[ 9973] = 64;
assign img[ 9974] = 54;
assign img[ 9975] = 64;
assign img[ 9976] = 64;
assign img[ 9977] = 64;
assign img[ 9978] = 56;
assign img[ 9979] = 64;
assign img[ 9980] = 56;
assign img[ 9981] = 64;
assign img[ 9982] = 58;
assign img[ 9983] = 64;
assign img[ 9984] = 64;
assign img[ 9985] = 86;
assign img[ 9986] = 81;
assign img[ 9987] = 84;
assign img[ 9988] = 90;
assign img[ 9989] = 87;
assign img[ 9990] = 96;
assign img[ 9991] = 88;
assign img[ 9992] = 96;
assign img[ 9993] = 98;
assign img[ 9994] = 98;
assign img[ 9995] = 100;
assign img[ 9996] = 101;
assign img[ 9997] = 101;
assign img[ 9998] = 102;
assign img[ 9999] = 110;
assign img[10000] = 97;
assign img[10001] = 98;
assign img[10002] = 98;
assign img[10003] = 97;
assign img[10004] = 102;
assign img[10005] = 97;
assign img[10006] = 101;
assign img[10007] = 104;
assign img[10008] = 104;
assign img[10009] = 97;
assign img[10010] = 102;
assign img[10011] = 100;
assign img[10012] = 101;
assign img[10013] = 93;
assign img[10014] = 97;
assign img[10015] = 95;
assign img[10016] = 104;
assign img[10017] = 97;
assign img[10018] = 106;
assign img[10019] = 101;
assign img[10020] = 104;
assign img[10021] = 100;
assign img[10022] = 101;
assign img[10023] = 103;
assign img[10024] = 98;
assign img[10025] = 97;
assign img[10026] = 97;
assign img[10027] = 101;
assign img[10028] = 97;
assign img[10029] = 97;
assign img[10030] = 101;
assign img[10031] = 104;
assign img[10032] = 104;
assign img[10033] = 97;
assign img[10034] = 101;
assign img[10035] = 104;
assign img[10036] = 96;
assign img[10037] = 97;
assign img[10038] = 100;
assign img[10039] = 100;
assign img[10040] = 100;
assign img[10041] = 101;
assign img[10042] = 100;
assign img[10043] = 96;
assign img[10044] = 101;
assign img[10045] = 96;
assign img[10046] = 109;
assign img[10047] = 101;
assign img[10048] = 97;
assign img[10049] = 109;
assign img[10050] = 101;
assign img[10051] = 97;
assign img[10052] = 104;
assign img[10053] = 96;
assign img[10054] = 77;
assign img[10055] = 83;
assign img[10056] = 81;
assign img[10057] = 81;
assign img[10058] = 73;
assign img[10059] = 78;
assign img[10060] = 76;
assign img[10061] = 73;
assign img[10062] = 80;
assign img[10063] = 84;
assign img[10064] = 72;
assign img[10065] = 72;
assign img[10066] = 68;
assign img[10067] = 72;
assign img[10068] = 77;
assign img[10069] = 70;
assign img[10070] = 73;
assign img[10071] = 76;
assign img[10072] = 74;
assign img[10073] = 80;
assign img[10074] = 71;
assign img[10075] = 69;
assign img[10076] = 76;
assign img[10077] = 76;
assign img[10078] = 76;
assign img[10079] = 73;
assign img[10080] = 70;
assign img[10081] = 86;
assign img[10082] = 77;
assign img[10083] = 76;
assign img[10084] = 76;
assign img[10085] = 76;
assign img[10086] = 66;
assign img[10087] = 72;
assign img[10088] = 78;
assign img[10089] = 72;
assign img[10090] = 68;
assign img[10091] = 70;
assign img[10092] = 70;
assign img[10093] = 68;
assign img[10094] = 70;
assign img[10095] = 78;
assign img[10096] = 68;
assign img[10097] = 66;
assign img[10098] = 71;
assign img[10099] = 70;
assign img[10100] = 76;
assign img[10101] = 70;
assign img[10102] = 71;
assign img[10103] = 64;
assign img[10104] = 66;
assign img[10105] = 68;
assign img[10106] = 72;
assign img[10107] = 71;
assign img[10108] = 64;
assign img[10109] = 76;
assign img[10110] = 68;
assign img[10111] = 68;
assign img[10112] = 69;
assign img[10113] = 64;
assign img[10114] = 64;
assign img[10115] = 56;
assign img[10116] = 64;
assign img[10117] = 64;
assign img[10118] = 65;
assign img[10119] = 64;
assign img[10120] = 66;
assign img[10121] = 73;
assign img[10122] = 81;
assign img[10123] = 83;
assign img[10124] = 74;
assign img[10125] = 83;
assign img[10126] = 77;
assign img[10127] = 77;
assign img[10128] = 81;
assign img[10129] = 75;
assign img[10130] = 79;
assign img[10131] = 77;
assign img[10132] = 81;
assign img[10133] = 81;
assign img[10134] = 81;
assign img[10135] = 81;
assign img[10136] = 81;
assign img[10137] = 82;
assign img[10138] = 88;
assign img[10139] = 84;
assign img[10140] = 84;
assign img[10141] = 73;
assign img[10142] = 83;
assign img[10143] = 83;
assign img[10144] = 80;
assign img[10145] = 81;
assign img[10146] = 74;
assign img[10147] = 73;
assign img[10148] = 81;
assign img[10149] = 79;
assign img[10150] = 73;
assign img[10151] = 75;
assign img[10152] = 73;
assign img[10153] = 78;
assign img[10154] = 81;
assign img[10155] = 70;
assign img[10156] = 84;
assign img[10157] = 69;
assign img[10158] = 81;
assign img[10159] = 77;
assign img[10160] = 81;
assign img[10161] = 83;
assign img[10162] = 80;
assign img[10163] = 81;
assign img[10164] = 80;
assign img[10165] = 73;
assign img[10166] = 74;
assign img[10167] = 77;
assign img[10168] = 77;
assign img[10169] = 76;
assign img[10170] = 77;
assign img[10171] = 83;
assign img[10172] = 80;
assign img[10173] = 83;
assign img[10174] = 84;
assign img[10175] = 80;
assign img[10176] = 81;
assign img[10177] = 81;
assign img[10178] = 75;
assign img[10179] = 85;
assign img[10180] = 69;
assign img[10181] = 77;
assign img[10182] = 70;
assign img[10183] = 65;
assign img[10184] = 57;
assign img[10185] = 56;
assign img[10186] = 54;
assign img[10187] = 57;
assign img[10188] = 60;
assign img[10189] = 57;
assign img[10190] = 58;
assign img[10191] = 53;
assign img[10192] = 45;
assign img[10193] = 57;
assign img[10194] = 53;
assign img[10195] = 58;
assign img[10196] = 54;
assign img[10197] = 50;
assign img[10198] = 51;
assign img[10199] = 45;
assign img[10200] = 48;
assign img[10201] = 54;
assign img[10202] = 60;
assign img[10203] = 52;
assign img[10204] = 51;
assign img[10205] = 64;
assign img[10206] = 54;
assign img[10207] = 52;
assign img[10208] = 45;
assign img[10209] = 50;
assign img[10210] = 50;
assign img[10211] = 56;
assign img[10212] = 51;
assign img[10213] = 54;
assign img[10214] = 50;
assign img[10215] = 55;
assign img[10216] = 53;
assign img[10217] = 51;
assign img[10218] = 49;
assign img[10219] = 57;
assign img[10220] = 53;
assign img[10221] = 50;
assign img[10222] = 52;
assign img[10223] = 54;
assign img[10224] = 49;
assign img[10225] = 48;
assign img[10226] = 60;
assign img[10227] = 55;
assign img[10228] = 53;
assign img[10229] = 53;
assign img[10230] = 55;
assign img[10231] = 49;
assign img[10232] = 47;
assign img[10233] = 49;
assign img[10234] = 52;
assign img[10235] = 50;
assign img[10236] = 53;
assign img[10237] = 53;
assign img[10238] = 52;
assign img[10239] = 53;
assign img[10240] = 33;
assign img[10241] = 45;
assign img[10242] = 48;
assign img[10243] = 52;
assign img[10244] = 46;
assign img[10245] = 54;
assign img[10246] = 54;
assign img[10247] = 64;
assign img[10248] = 64;
assign img[10249] = 68;
assign img[10250] = 71;
assign img[10251] = 71;
assign img[10252] = 71;
assign img[10253] = 72;
assign img[10254] = 69;
assign img[10255] = 71;
assign img[10256] = 76;
assign img[10257] = 65;
assign img[10258] = 75;
assign img[10259] = 64;
assign img[10260] = 72;
assign img[10261] = 79;
assign img[10262] = 65;
assign img[10263] = 68;
assign img[10264] = 64;
assign img[10265] = 64;
assign img[10266] = 66;
assign img[10267] = 66;
assign img[10268] = 70;
assign img[10269] = 66;
assign img[10270] = 67;
assign img[10271] = 75;
assign img[10272] = 68;
assign img[10273] = 68;
assign img[10274] = 66;
assign img[10275] = 73;
assign img[10276] = 70;
assign img[10277] = 70;
assign img[10278] = 68;
assign img[10279] = 70;
assign img[10280] = 68;
assign img[10281] = 64;
assign img[10282] = 66;
assign img[10283] = 66;
assign img[10284] = 68;
assign img[10285] = 73;
assign img[10286] = 66;
assign img[10287] = 72;
assign img[10288] = 71;
assign img[10289] = 76;
assign img[10290] = 70;
assign img[10291] = 70;
assign img[10292] = 70;
assign img[10293] = 68;
assign img[10294] = 64;
assign img[10295] = 66;
assign img[10296] = 70;
assign img[10297] = 74;
assign img[10298] = 68;
assign img[10299] = 74;
assign img[10300] = 69;
assign img[10301] = 64;
assign img[10302] = 78;
assign img[10303] = 76;
assign img[10304] = 68;
assign img[10305] = 68;
assign img[10306] = 68;
assign img[10307] = 64;
assign img[10308] = 64;
assign img[10309] = 65;
assign img[10310] = 67;
assign img[10311] = 64;
assign img[10312] = 64;
assign img[10313] = 47;
assign img[10314] = 46;
assign img[10315] = 46;
assign img[10316] = 42;
assign img[10317] = 46;
assign img[10318] = 47;
assign img[10319] = 44;
assign img[10320] = 44;
assign img[10321] = 42;
assign img[10322] = 38;
assign img[10323] = 42;
assign img[10324] = 45;
assign img[10325] = 41;
assign img[10326] = 48;
assign img[10327] = 39;
assign img[10328] = 44;
assign img[10329] = 37;
assign img[10330] = 40;
assign img[10331] = 39;
assign img[10332] = 38;
assign img[10333] = 38;
assign img[10334] = 38;
assign img[10335] = 36;
assign img[10336] = 38;
assign img[10337] = 42;
assign img[10338] = 44;
assign img[10339] = 38;
assign img[10340] = 38;
assign img[10341] = 36;
assign img[10342] = 40;
assign img[10343] = 33;
assign img[10344] = 38;
assign img[10345] = 39;
assign img[10346] = 44;
assign img[10347] = 44;
assign img[10348] = 38;
assign img[10349] = 38;
assign img[10350] = 38;
assign img[10351] = 44;
assign img[10352] = 32;
assign img[10353] = 34;
assign img[10354] = 38;
assign img[10355] = 40;
assign img[10356] = 40;
assign img[10357] = 36;
assign img[10358] = 36;
assign img[10359] = 36;
assign img[10360] = 36;
assign img[10361] = 36;
assign img[10362] = 38;
assign img[10363] = 38;
assign img[10364] = 38;
assign img[10365] = 44;
assign img[10366] = 38;
assign img[10367] = 42;
assign img[10368] = 38;
assign img[10369] = 54;
assign img[10370] = 64;
assign img[10371] = 50;
assign img[10372] = 54;
assign img[10373] = 51;
assign img[10374] = 58;
assign img[10375] = 70;
assign img[10376] = 65;
assign img[10377] = 69;
assign img[10378] = 76;
assign img[10379] = 79;
assign img[10380] = 76;
assign img[10381] = 72;
assign img[10382] = 78;
assign img[10383] = 77;
assign img[10384] = 70;
assign img[10385] = 78;
assign img[10386] = 84;
assign img[10387] = 72;
assign img[10388] = 78;
assign img[10389] = 78;
assign img[10390] = 79;
assign img[10391] = 78;
assign img[10392] = 76;
assign img[10393] = 80;
assign img[10394] = 86;
assign img[10395] = 78;
assign img[10396] = 79;
assign img[10397] = 71;
assign img[10398] = 76;
assign img[10399] = 86;
assign img[10400] = 78;
assign img[10401] = 86;
assign img[10402] = 86;
assign img[10403] = 76;
assign img[10404] = 70;
assign img[10405] = 79;
assign img[10406] = 80;
assign img[10407] = 77;
assign img[10408] = 79;
assign img[10409] = 80;
assign img[10410] = 78;
assign img[10411] = 79;
assign img[10412] = 71;
assign img[10413] = 78;
assign img[10414] = 78;
assign img[10415] = 72;
assign img[10416] = 80;
assign img[10417] = 86;
assign img[10418] = 78;
assign img[10419] = 79;
assign img[10420] = 78;
assign img[10421] = 80;
assign img[10422] = 78;
assign img[10423] = 71;
assign img[10424] = 72;
assign img[10425] = 76;
assign img[10426] = 72;
assign img[10427] = 71;
assign img[10428] = 72;
assign img[10429] = 72;
assign img[10430] = 75;
assign img[10431] = 76;
assign img[10432] = 70;
assign img[10433] = 73;
assign img[10434] = 72;
assign img[10435] = 76;
assign img[10436] = 70;
assign img[10437] = 72;
assign img[10438] = 69;
assign img[10439] = 68;
assign img[10440] = 64;
assign img[10441] = 64;
assign img[10442] = 54;
assign img[10443] = 47;
assign img[10444] = 46;
assign img[10445] = 46;
assign img[10446] = 47;
assign img[10447] = 44;
assign img[10448] = 52;
assign img[10449] = 51;
assign img[10450] = 48;
assign img[10451] = 48;
assign img[10452] = 54;
assign img[10453] = 48;
assign img[10454] = 52;
assign img[10455] = 48;
assign img[10456] = 48;
assign img[10457] = 44;
assign img[10458] = 45;
assign img[10459] = 46;
assign img[10460] = 46;
assign img[10461] = 50;
assign img[10462] = 52;
assign img[10463] = 48;
assign img[10464] = 42;
assign img[10465] = 44;
assign img[10466] = 52;
assign img[10467] = 52;
assign img[10468] = 47;
assign img[10469] = 44;
assign img[10470] = 48;
assign img[10471] = 50;
assign img[10472] = 47;
assign img[10473] = 40;
assign img[10474] = 45;
assign img[10475] = 52;
assign img[10476] = 51;
assign img[10477] = 49;
assign img[10478] = 44;
assign img[10479] = 48;
assign img[10480] = 44;
assign img[10481] = 47;
assign img[10482] = 44;
assign img[10483] = 40;
assign img[10484] = 40;
assign img[10485] = 41;
assign img[10486] = 44;
assign img[10487] = 40;
assign img[10488] = 44;
assign img[10489] = 44;
assign img[10490] = 40;
assign img[10491] = 44;
assign img[10492] = 44;
assign img[10493] = 46;
assign img[10494] = 52;
assign img[10495] = 43;
assign img[10496] = 44;
assign img[10497] = 31;
assign img[10498] = 30;
assign img[10499] = 29;
assign img[10500] = 28;
assign img[10501] = 30;
assign img[10502] = 31;
assign img[10503] = 38;
assign img[10504] = 47;
assign img[10505] = 44;
assign img[10506] = 48;
assign img[10507] = 48;
assign img[10508] = 46;
assign img[10509] = 47;
assign img[10510] = 55;
assign img[10511] = 48;
assign img[10512] = 48;
assign img[10513] = 46;
assign img[10514] = 48;
assign img[10515] = 46;
assign img[10516] = 43;
assign img[10517] = 42;
assign img[10518] = 48;
assign img[10519] = 46;
assign img[10520] = 46;
assign img[10521] = 46;
assign img[10522] = 41;
assign img[10523] = 46;
assign img[10524] = 46;
assign img[10525] = 47;
assign img[10526] = 48;
assign img[10527] = 44;
assign img[10528] = 47;
assign img[10529] = 52;
assign img[10530] = 47;
assign img[10531] = 46;
assign img[10532] = 45;
assign img[10533] = 48;
assign img[10534] = 45;
assign img[10535] = 47;
assign img[10536] = 47;
assign img[10537] = 52;
assign img[10538] = 47;
assign img[10539] = 52;
assign img[10540] = 46;
assign img[10541] = 47;
assign img[10542] = 49;
assign img[10543] = 46;
assign img[10544] = 47;
assign img[10545] = 54;
assign img[10546] = 43;
assign img[10547] = 52;
assign img[10548] = 54;
assign img[10549] = 47;
assign img[10550] = 40;
assign img[10551] = 51;
assign img[10552] = 42;
assign img[10553] = 46;
assign img[10554] = 55;
assign img[10555] = 53;
assign img[10556] = 47;
assign img[10557] = 43;
assign img[10558] = 43;
assign img[10559] = 48;
assign img[10560] = 45;
assign img[10561] = 48;
assign img[10562] = 41;
assign img[10563] = 50;
assign img[10564] = 47;
assign img[10565] = 46;
assign img[10566] = 41;
assign img[10567] = 37;
assign img[10568] = 40;
assign img[10569] = 39;
assign img[10570] = 33;
assign img[10571] = 25;
assign img[10572] = 28;
assign img[10573] = 28;
assign img[10574] = 29;
assign img[10575] = 29;
assign img[10576] = 25;
assign img[10577] = 26;
assign img[10578] = 22;
assign img[10579] = 26;
assign img[10580] = 26;
assign img[10581] = 28;
assign img[10582] = 29;
assign img[10583] = 24;
assign img[10584] = 19;
assign img[10585] = 21;
assign img[10586] = 26;
assign img[10587] = 23;
assign img[10588] = 22;
assign img[10589] = 20;
assign img[10590] = 24;
assign img[10591] = 20;
assign img[10592] = 18;
assign img[10593] = 24;
assign img[10594] = 26;
assign img[10595] = 22;
assign img[10596] = 16;
assign img[10597] = 18;
assign img[10598] = 16;
assign img[10599] = 20;
assign img[10600] = 20;
assign img[10601] = 26;
assign img[10602] = 28;
assign img[10603] = 21;
assign img[10604] = 21;
assign img[10605] = 17;
assign img[10606] = 22;
assign img[10607] = 21;
assign img[10608] = 24;
assign img[10609] = 18;
assign img[10610] = 21;
assign img[10611] = 18;
assign img[10612] = 16;
assign img[10613] = 16;
assign img[10614] = 20;
assign img[10615] = 19;
assign img[10616] = 22;
assign img[10617] = 21;
assign img[10618] = 17;
assign img[10619] = 16;
assign img[10620] = 18;
assign img[10621] = 16;
assign img[10622] = 24;
assign img[10623] = 15;
assign img[10624] = 18;
assign img[10625] = 68;
assign img[10626] = 69;
assign img[10627] = 66;
assign img[10628] = 65;
assign img[10629] = 65;
assign img[10630] = 69;
assign img[10631] = 82;
assign img[10632] = 86;
assign img[10633] = 92;
assign img[10634] = 88;
assign img[10635] = 88;
assign img[10636] = 94;
assign img[10637] = 88;
assign img[10638] = 86;
assign img[10639] = 99;
assign img[10640] = 92;
assign img[10641] = 88;
assign img[10642] = 90;
assign img[10643] = 86;
assign img[10644] = 87;
assign img[10645] = 88;
assign img[10646] = 86;
assign img[10647] = 92;
assign img[10648] = 88;
assign img[10649] = 86;
assign img[10650] = 95;
assign img[10651] = 90;
assign img[10652] = 86;
assign img[10653] = 86;
assign img[10654] = 86;
assign img[10655] = 88;
assign img[10656] = 92;
assign img[10657] = 87;
assign img[10658] = 90;
assign img[10659] = 88;
assign img[10660] = 100;
assign img[10661] = 87;
assign img[10662] = 94;
assign img[10663] = 88;
assign img[10664] = 94;
assign img[10665] = 84;
assign img[10666] = 96;
assign img[10667] = 98;
assign img[10668] = 87;
assign img[10669] = 86;
assign img[10670] = 87;
assign img[10671] = 91;
assign img[10672] = 87;
assign img[10673] = 87;
assign img[10674] = 86;
assign img[10675] = 86;
assign img[10676] = 90;
assign img[10677] = 86;
assign img[10678] = 86;
assign img[10679] = 96;
assign img[10680] = 88;
assign img[10681] = 94;
assign img[10682] = 92;
assign img[10683] = 87;
assign img[10684] = 90;
assign img[10685] = 84;
assign img[10686] = 80;
assign img[10687] = 92;
assign img[10688] = 81;
assign img[10689] = 82;
assign img[10690] = 85;
assign img[10691] = 84;
assign img[10692] = 81;
assign img[10693] = 86;
assign img[10694] = 92;
assign img[10695] = 84;
assign img[10696] = 80;
assign img[10697] = 73;
assign img[10698] = 70;
assign img[10699] = 65;
assign img[10700] = 74;
assign img[10701] = 65;
assign img[10702] = 67;
assign img[10703] = 64;
assign img[10704] = 64;
assign img[10705] = 64;
assign img[10706] = 65;
assign img[10707] = 69;
assign img[10708] = 64;
assign img[10709] = 64;
assign img[10710] = 65;
assign img[10711] = 64;
assign img[10712] = 54;
assign img[10713] = 64;
assign img[10714] = 52;
assign img[10715] = 64;
assign img[10716] = 64;
assign img[10717] = 56;
assign img[10718] = 64;
assign img[10719] = 64;
assign img[10720] = 64;
assign img[10721] = 64;
assign img[10722] = 54;
assign img[10723] = 64;
assign img[10724] = 64;
assign img[10725] = 64;
assign img[10726] = 64;
assign img[10727] = 64;
assign img[10728] = 64;
assign img[10729] = 65;
assign img[10730] = 64;
assign img[10731] = 64;
assign img[10732] = 55;
assign img[10733] = 64;
assign img[10734] = 65;
assign img[10735] = 53;
assign img[10736] = 64;
assign img[10737] = 64;
assign img[10738] = 58;
assign img[10739] = 64;
assign img[10740] = 52;
assign img[10741] = 64;
assign img[10742] = 53;
assign img[10743] = 51;
assign img[10744] = 48;
assign img[10745] = 52;
assign img[10746] = 64;
assign img[10747] = 64;
assign img[10748] = 53;
assign img[10749] = 56;
assign img[10750] = 54;
assign img[10751] = 64;
assign img[10752] = 46;
assign img[10753] = 68;
assign img[10754] = 68;
assign img[10755] = 66;
assign img[10756] = 64;
assign img[10757] = 65;
assign img[10758] = 68;
assign img[10759] = 73;
assign img[10760] = 77;
assign img[10761] = 78;
assign img[10762] = 84;
assign img[10763] = 87;
assign img[10764] = 94;
assign img[10765] = 79;
assign img[10766] = 86;
assign img[10767] = 82;
assign img[10768] = 80;
assign img[10769] = 92;
assign img[10770] = 86;
assign img[10771] = 86;
assign img[10772] = 86;
assign img[10773] = 87;
assign img[10774] = 84;
assign img[10775] = 86;
assign img[10776] = 87;
assign img[10777] = 86;
assign img[10778] = 86;
assign img[10779] = 85;
assign img[10780] = 84;
assign img[10781] = 78;
assign img[10782] = 92;
assign img[10783] = 86;
assign img[10784] = 84;
assign img[10785] = 88;
assign img[10786] = 80;
assign img[10787] = 96;
assign img[10788] = 81;
assign img[10789] = 88;
assign img[10790] = 86;
assign img[10791] = 80;
assign img[10792] = 84;
assign img[10793] = 88;
assign img[10794] = 87;
assign img[10795] = 86;
assign img[10796] = 79;
assign img[10797] = 78;
assign img[10798] = 84;
assign img[10799] = 86;
assign img[10800] = 94;
assign img[10801] = 80;
assign img[10802] = 86;
assign img[10803] = 86;
assign img[10804] = 84;
assign img[10805] = 86;
assign img[10806] = 82;
assign img[10807] = 87;
assign img[10808] = 86;
assign img[10809] = 84;
assign img[10810] = 86;
assign img[10811] = 86;
assign img[10812] = 82;
assign img[10813] = 85;
assign img[10814] = 80;
assign img[10815] = 80;
assign img[10816] = 77;
assign img[10817] = 79;
assign img[10818] = 84;
assign img[10819] = 84;
assign img[10820] = 79;
assign img[10821] = 88;
assign img[10822] = 84;
assign img[10823] = 79;
assign img[10824] = 78;
assign img[10825] = 79;
assign img[10826] = 72;
assign img[10827] = 65;
assign img[10828] = 64;
assign img[10829] = 57;
assign img[10830] = 64;
assign img[10831] = 65;
assign img[10832] = 64;
assign img[10833] = 64;
assign img[10834] = 64;
assign img[10835] = 64;
assign img[10836] = 65;
assign img[10837] = 64;
assign img[10838] = 57;
assign img[10839] = 64;
assign img[10840] = 64;
assign img[10841] = 65;
assign img[10842] = 64;
assign img[10843] = 58;
assign img[10844] = 64;
assign img[10845] = 57;
assign img[10846] = 64;
assign img[10847] = 57;
assign img[10848] = 53;
assign img[10849] = 53;
assign img[10850] = 64;
assign img[10851] = 57;
assign img[10852] = 64;
assign img[10853] = 57;
assign img[10854] = 53;
assign img[10855] = 52;
assign img[10856] = 54;
assign img[10857] = 52;
assign img[10858] = 48;
assign img[10859] = 55;
assign img[10860] = 64;
assign img[10861] = 52;
assign img[10862] = 56;
assign img[10863] = 53;
assign img[10864] = 56;
assign img[10865] = 51;
assign img[10866] = 52;
assign img[10867] = 55;
assign img[10868] = 56;
assign img[10869] = 64;
assign img[10870] = 45;
assign img[10871] = 52;
assign img[10872] = 64;
assign img[10873] = 52;
assign img[10874] = 56;
assign img[10875] = 52;
assign img[10876] = 52;
assign img[10877] = 57;
assign img[10878] = 54;
assign img[10879] = 52;
assign img[10880] = 51;
assign img[10881] = 64;
assign img[10882] = 51;
assign img[10883] = 53;
assign img[10884] = 64;
assign img[10885] = 56;
assign img[10886] = 76;
assign img[10887] = 68;
assign img[10888] = 72;
assign img[10889] = 72;
assign img[10890] = 70;
assign img[10891] = 72;
assign img[10892] = 79;
assign img[10893] = 72;
assign img[10894] = 70;
assign img[10895] = 78;
assign img[10896] = 70;
assign img[10897] = 72;
assign img[10898] = 79;
assign img[10899] = 79;
assign img[10900] = 76;
assign img[10901] = 72;
assign img[10902] = 72;
assign img[10903] = 71;
assign img[10904] = 76;
assign img[10905] = 79;
assign img[10906] = 80;
assign img[10907] = 78;
assign img[10908] = 76;
assign img[10909] = 80;
assign img[10910] = 78;
assign img[10911] = 78;
assign img[10912] = 72;
assign img[10913] = 82;
assign img[10914] = 72;
assign img[10915] = 78;
assign img[10916] = 71;
assign img[10917] = 72;
assign img[10918] = 72;
assign img[10919] = 80;
assign img[10920] = 79;
assign img[10921] = 75;
assign img[10922] = 78;
assign img[10923] = 78;
assign img[10924] = 72;
assign img[10925] = 78;
assign img[10926] = 86;
assign img[10927] = 72;
assign img[10928] = 69;
assign img[10929] = 75;
assign img[10930] = 79;
assign img[10931] = 86;
assign img[10932] = 73;
assign img[10933] = 72;
assign img[10934] = 78;
assign img[10935] = 78;
assign img[10936] = 72;
assign img[10937] = 76;
assign img[10938] = 77;
assign img[10939] = 72;
assign img[10940] = 71;
assign img[10941] = 72;
assign img[10942] = 76;
assign img[10943] = 72;
assign img[10944] = 72;
assign img[10945] = 69;
assign img[10946] = 72;
assign img[10947] = 76;
assign img[10948] = 69;
assign img[10949] = 75;
assign img[10950] = 72;
assign img[10951] = 65;
assign img[10952] = 72;
assign img[10953] = 68;
assign img[10954] = 64;
assign img[10955] = 70;
assign img[10956] = 50;
assign img[10957] = 49;
assign img[10958] = 46;
assign img[10959] = 46;
assign img[10960] = 47;
assign img[10961] = 47;
assign img[10962] = 46;
assign img[10963] = 52;
assign img[10964] = 48;
assign img[10965] = 47;
assign img[10966] = 50;
assign img[10967] = 46;
assign img[10968] = 41;
assign img[10969] = 47;
assign img[10970] = 52;
assign img[10971] = 52;
assign img[10972] = 46;
assign img[10973] = 41;
assign img[10974] = 52;
assign img[10975] = 45;
assign img[10976] = 42;
assign img[10977] = 49;
assign img[10978] = 45;
assign img[10979] = 64;
assign img[10980] = 42;
assign img[10981] = 48;
assign img[10982] = 49;
assign img[10983] = 50;
assign img[10984] = 45;
assign img[10985] = 48;
assign img[10986] = 49;
assign img[10987] = 44;
assign img[10988] = 45;
assign img[10989] = 44;
assign img[10990] = 46;
assign img[10991] = 44;
assign img[10992] = 40;
assign img[10993] = 46;
assign img[10994] = 44;
assign img[10995] = 40;
assign img[10996] = 44;
assign img[10997] = 41;
assign img[10998] = 43;
assign img[10999] = 42;
assign img[11000] = 41;
assign img[11001] = 44;
assign img[11002] = 45;
assign img[11003] = 45;
assign img[11004] = 41;
assign img[11005] = 49;
assign img[11006] = 45;
assign img[11007] = 40;
assign img[11008] = 46;
assign img[11009] = 44;
assign img[11010] = 44;
assign img[11011] = 44;
assign img[11012] = 44;
assign img[11013] = 52;
assign img[11014] = 48;
assign img[11015] = 53;
assign img[11016] = 64;
assign img[11017] = 64;
assign img[11018] = 65;
assign img[11019] = 64;
assign img[11020] = 64;
assign img[11021] = 67;
assign img[11022] = 68;
assign img[11023] = 64;
assign img[11024] = 64;
assign img[11025] = 64;
assign img[11026] = 64;
assign img[11027] = 64;
assign img[11028] = 64;
assign img[11029] = 64;
assign img[11030] = 64;
assign img[11031] = 64;
assign img[11032] = 65;
assign img[11033] = 68;
assign img[11034] = 64;
assign img[11035] = 66;
assign img[11036] = 64;
assign img[11037] = 69;
assign img[11038] = 69;
assign img[11039] = 64;
assign img[11040] = 64;
assign img[11041] = 67;
assign img[11042] = 68;
assign img[11043] = 64;
assign img[11044] = 65;
assign img[11045] = 64;
assign img[11046] = 70;
assign img[11047] = 64;
assign img[11048] = 65;
assign img[11049] = 65;
assign img[11050] = 65;
assign img[11051] = 64;
assign img[11052] = 69;
assign img[11053] = 64;
assign img[11054] = 66;
assign img[11055] = 64;
assign img[11056] = 65;
assign img[11057] = 65;
assign img[11058] = 64;
assign img[11059] = 65;
assign img[11060] = 66;
assign img[11061] = 64;
assign img[11062] = 66;
assign img[11063] = 64;
assign img[11064] = 64;
assign img[11065] = 64;
assign img[11066] = 64;
assign img[11067] = 64;
assign img[11068] = 64;
assign img[11069] = 65;
assign img[11070] = 64;
assign img[11071] = 66;
assign img[11072] = 65;
assign img[11073] = 64;
assign img[11074] = 67;
assign img[11075] = 64;
assign img[11076] = 65;
assign img[11077] = 69;
assign img[11078] = 65;
assign img[11079] = 64;
assign img[11080] = 64;
assign img[11081] = 68;
assign img[11082] = 64;
assign img[11083] = 53;
assign img[11084] = 52;
assign img[11085] = 42;
assign img[11086] = 45;
assign img[11087] = 40;
assign img[11088] = 36;
assign img[11089] = 47;
assign img[11090] = 46;
assign img[11091] = 46;
assign img[11092] = 41;
assign img[11093] = 44;
assign img[11094] = 37;
assign img[11095] = 38;
assign img[11096] = 40;
assign img[11097] = 39;
assign img[11098] = 41;
assign img[11099] = 41;
assign img[11100] = 41;
assign img[11101] = 39;
assign img[11102] = 38;
assign img[11103] = 41;
assign img[11104] = 37;
assign img[11105] = 41;
assign img[11106] = 38;
assign img[11107] = 38;
assign img[11108] = 37;
assign img[11109] = 35;
assign img[11110] = 41;
assign img[11111] = 34;
assign img[11112] = 36;
assign img[11113] = 36;
assign img[11114] = 40;
assign img[11115] = 36;
assign img[11116] = 34;
assign img[11117] = 38;
assign img[11118] = 40;
assign img[11119] = 37;
assign img[11120] = 39;
assign img[11121] = 37;
assign img[11122] = 42;
assign img[11123] = 39;
assign img[11124] = 32;
assign img[11125] = 35;
assign img[11126] = 36;
assign img[11127] = 34;
assign img[11128] = 30;
assign img[11129] = 36;
assign img[11130] = 36;
assign img[11131] = 38;
assign img[11132] = 38;
assign img[11133] = 34;
assign img[11134] = 39;
assign img[11135] = 33;
assign img[11136] = 32;
assign img[11137] = 53;
assign img[11138] = 64;
assign img[11139] = 52;
assign img[11140] = 56;
assign img[11141] = 64;
assign img[11142] = 65;
assign img[11143] = 66;
assign img[11144] = 72;
assign img[11145] = 69;
assign img[11146] = 79;
assign img[11147] = 70;
assign img[11148] = 77;
assign img[11149] = 73;
assign img[11150] = 74;
assign img[11151] = 73;
assign img[11152] = 69;
assign img[11153] = 73;
assign img[11154] = 74;
assign img[11155] = 78;
assign img[11156] = 72;
assign img[11157] = 72;
assign img[11158] = 73;
assign img[11159] = 77;
assign img[11160] = 73;
assign img[11161] = 73;
assign img[11162] = 79;
assign img[11163] = 73;
assign img[11164] = 74;
assign img[11165] = 77;
assign img[11166] = 71;
assign img[11167] = 72;
assign img[11168] = 73;
assign img[11169] = 77;
assign img[11170] = 77;
assign img[11171] = 70;
assign img[11172] = 76;
assign img[11173] = 88;
assign img[11174] = 77;
assign img[11175] = 73;
assign img[11176] = 74;
assign img[11177] = 80;
assign img[11178] = 71;
assign img[11179] = 73;
assign img[11180] = 73;
assign img[11181] = 74;
assign img[11182] = 77;
assign img[11183] = 77;
assign img[11184] = 77;
assign img[11185] = 81;
assign img[11186] = 77;
assign img[11187] = 78;
assign img[11188] = 77;
assign img[11189] = 77;
assign img[11190] = 80;
assign img[11191] = 73;
assign img[11192] = 72;
assign img[11193] = 74;
assign img[11194] = 72;
assign img[11195] = 73;
assign img[11196] = 77;
assign img[11197] = 78;
assign img[11198] = 77;
assign img[11199] = 73;
assign img[11200] = 74;
assign img[11201] = 79;
assign img[11202] = 72;
assign img[11203] = 80;
assign img[11204] = 66;
assign img[11205] = 79;
assign img[11206] = 77;
assign img[11207] = 77;
assign img[11208] = 73;
assign img[11209] = 69;
assign img[11210] = 73;
assign img[11211] = 73;
assign img[11212] = 65;
assign img[11213] = 65;
assign img[11214] = 53;
assign img[11215] = 57;
assign img[11216] = 51;
assign img[11217] = 54;
assign img[11218] = 47;
assign img[11219] = 56;
assign img[11220] = 53;
assign img[11221] = 49;
assign img[11222] = 50;
assign img[11223] = 52;
assign img[11224] = 52;
assign img[11225] = 46;
assign img[11226] = 53;
assign img[11227] = 47;
assign img[11228] = 47;
assign img[11229] = 44;
assign img[11230] = 46;
assign img[11231] = 44;
assign img[11232] = 46;
assign img[11233] = 52;
assign img[11234] = 45;
assign img[11235] = 41;
assign img[11236] = 44;
assign img[11237] = 45;
assign img[11238] = 45;
assign img[11239] = 45;
assign img[11240] = 44;
assign img[11241] = 44;
assign img[11242] = 48;
assign img[11243] = 44;
assign img[11244] = 46;
assign img[11245] = 41;
assign img[11246] = 47;
assign img[11247] = 52;
assign img[11248] = 42;
assign img[11249] = 45;
assign img[11250] = 45;
assign img[11251] = 40;
assign img[11252] = 44;
assign img[11253] = 44;
assign img[11254] = 48;
assign img[11255] = 44;
assign img[11256] = 42;
assign img[11257] = 48;
assign img[11258] = 44;
assign img[11259] = 46;
assign img[11260] = 48;
assign img[11261] = 47;
assign img[11262] = 45;
assign img[11263] = 45;
assign img[11264] = 44;
assign img[11265] = 47;
assign img[11266] = 47;
assign img[11267] = 45;
assign img[11268] = 46;
assign img[11269] = 54;
assign img[11270] = 64;
assign img[11271] = 53;
assign img[11272] = 65;
assign img[11273] = 64;
assign img[11274] = 64;
assign img[11275] = 68;
assign img[11276] = 65;
assign img[11277] = 65;
assign img[11278] = 77;
assign img[11279] = 73;
assign img[11280] = 53;
assign img[11281] = 69;
assign img[11282] = 72;
assign img[11283] = 67;
assign img[11284] = 65;
assign img[11285] = 66;
assign img[11286] = 73;
assign img[11287] = 65;
assign img[11288] = 64;
assign img[11289] = 73;
assign img[11290] = 71;
assign img[11291] = 68;
assign img[11292] = 69;
assign img[11293] = 65;
assign img[11294] = 66;
assign img[11295] = 72;
assign img[11296] = 67;
assign img[11297] = 69;
assign img[11298] = 74;
assign img[11299] = 64;
assign img[11300] = 67;
assign img[11301] = 71;
assign img[11302] = 64;
assign img[11303] = 69;
assign img[11304] = 66;
assign img[11305] = 72;
assign img[11306] = 69;
assign img[11307] = 64;
assign img[11308] = 65;
assign img[11309] = 68;
assign img[11310] = 66;
assign img[11311] = 70;
assign img[11312] = 69;
assign img[11313] = 72;
assign img[11314] = 66;
assign img[11315] = 73;
assign img[11316] = 65;
assign img[11317] = 64;
assign img[11318] = 65;
assign img[11319] = 65;
assign img[11320] = 68;
assign img[11321] = 69;
assign img[11322] = 66;
assign img[11323] = 71;
assign img[11324] = 69;
assign img[11325] = 65;
assign img[11326] = 69;
assign img[11327] = 66;
assign img[11328] = 70;
assign img[11329] = 65;
assign img[11330] = 66;
assign img[11331] = 66;
assign img[11332] = 65;
assign img[11333] = 72;
assign img[11334] = 66;
assign img[11335] = 67;
assign img[11336] = 66;
assign img[11337] = 70;
assign img[11338] = 65;
assign img[11339] = 64;
assign img[11340] = 58;
assign img[11341] = 52;
assign img[11342] = 52;
assign img[11343] = 48;
assign img[11344] = 44;
assign img[11345] = 45;
assign img[11346] = 48;
assign img[11347] = 45;
assign img[11348] = 42;
assign img[11349] = 45;
assign img[11350] = 51;
assign img[11351] = 49;
assign img[11352] = 46;
assign img[11353] = 44;
assign img[11354] = 48;
assign img[11355] = 39;
assign img[11356] = 45;
assign img[11357] = 44;
assign img[11358] = 39;
assign img[11359] = 44;
assign img[11360] = 39;
assign img[11361] = 42;
assign img[11362] = 44;
assign img[11363] = 41;
assign img[11364] = 44;
assign img[11365] = 45;
assign img[11366] = 39;
assign img[11367] = 41;
assign img[11368] = 46;
assign img[11369] = 45;
assign img[11370] = 45;
assign img[11371] = 41;
assign img[11372] = 39;
assign img[11373] = 41;
assign img[11374] = 38;
assign img[11375] = 44;
assign img[11376] = 37;
assign img[11377] = 34;
assign img[11378] = 41;
assign img[11379] = 38;
assign img[11380] = 41;
assign img[11381] = 35;
assign img[11382] = 37;
assign img[11383] = 37;
assign img[11384] = 39;
assign img[11385] = 40;
assign img[11386] = 41;
assign img[11387] = 38;
assign img[11388] = 34;
assign img[11389] = 37;
assign img[11390] = 39;
assign img[11391] = 37;
assign img[11392] = 44;
assign img[11393] = 29;
assign img[11394] = 33;
assign img[11395] = 30;
assign img[11396] = 34;
assign img[11397] = 33;
assign img[11398] = 45;
assign img[11399] = 48;
assign img[11400] = 44;
assign img[11401] = 48;
assign img[11402] = 49;
assign img[11403] = 56;
assign img[11404] = 44;
assign img[11405] = 52;
assign img[11406] = 45;
assign img[11407] = 52;
assign img[11408] = 50;
assign img[11409] = 49;
assign img[11410] = 52;
assign img[11411] = 48;
assign img[11412] = 50;
assign img[11413] = 46;
assign img[11414] = 52;
assign img[11415] = 46;
assign img[11416] = 44;
assign img[11417] = 44;
assign img[11418] = 47;
assign img[11419] = 44;
assign img[11420] = 44;
assign img[11421] = 52;
assign img[11422] = 46;
assign img[11423] = 56;
assign img[11424] = 53;
assign img[11425] = 51;
assign img[11426] = 48;
assign img[11427] = 48;
assign img[11428] = 49;
assign img[11429] = 52;
assign img[11430] = 52;
assign img[11431] = 43;
assign img[11432] = 48;
assign img[11433] = 47;
assign img[11434] = 53;
assign img[11435] = 51;
assign img[11436] = 52;
assign img[11437] = 41;
assign img[11438] = 52;
assign img[11439] = 46;
assign img[11440] = 46;
assign img[11441] = 48;
assign img[11442] = 45;
assign img[11443] = 52;
assign img[11444] = 52;
assign img[11445] = 50;
assign img[11446] = 50;
assign img[11447] = 51;
assign img[11448] = 48;
assign img[11449] = 47;
assign img[11450] = 48;
assign img[11451] = 46;
assign img[11452] = 42;
assign img[11453] = 50;
assign img[11454] = 52;
assign img[11455] = 45;
assign img[11456] = 46;
assign img[11457] = 52;
assign img[11458] = 48;
assign img[11459] = 46;
assign img[11460] = 45;
assign img[11461] = 48;
assign img[11462] = 44;
assign img[11463] = 43;
assign img[11464] = 46;
assign img[11465] = 48;
assign img[11466] = 49;
assign img[11467] = 48;
assign img[11468] = 37;
assign img[11469] = 44;
assign img[11470] = 34;
assign img[11471] = 35;
assign img[11472] = 28;
assign img[11473] = 32;
assign img[11474] = 29;
assign img[11475] = 32;
assign img[11476] = 33;
assign img[11477] = 27;
assign img[11478] = 25;
assign img[11479] = 24;
assign img[11480] = 20;
assign img[11481] = 24;
assign img[11482] = 28;
assign img[11483] = 27;
assign img[11484] = 26;
assign img[11485] = 26;
assign img[11486] = 32;
assign img[11487] = 32;
assign img[11488] = 27;
assign img[11489] = 28;
assign img[11490] = 24;
assign img[11491] = 26;
assign img[11492] = 26;
assign img[11493] = 24;
assign img[11494] = 32;
assign img[11495] = 24;
assign img[11496] = 29;
assign img[11497] = 28;
assign img[11498] = 23;
assign img[11499] = 28;
assign img[11500] = 25;
assign img[11501] = 28;
assign img[11502] = 21;
assign img[11503] = 27;
assign img[11504] = 22;
assign img[11505] = 22;
assign img[11506] = 24;
assign img[11507] = 24;
assign img[11508] = 25;
assign img[11509] = 23;
assign img[11510] = 22;
assign img[11511] = 29;
assign img[11512] = 18;
assign img[11513] = 22;
assign img[11514] = 27;
assign img[11515] = 26;
assign img[11516] = 23;
assign img[11517] = 28;
assign img[11518] = 23;
assign img[11519] = 27;
assign img[11520] = 25;
assign img[11521] = 67;
assign img[11522] = 64;
assign img[11523] = 64;
assign img[11524] = 64;
assign img[11525] = 64;
assign img[11526] = 77;
assign img[11527] = 72;
assign img[11528] = 72;
assign img[11529] = 75;
assign img[11530] = 77;
assign img[11531] = 80;
assign img[11532] = 78;
assign img[11533] = 81;
assign img[11534] = 74;
assign img[11535] = 78;
assign img[11536] = 77;
assign img[11537] = 78;
assign img[11538] = 77;
assign img[11539] = 76;
assign img[11540] = 82;
assign img[11541] = 79;
assign img[11542] = 73;
assign img[11543] = 80;
assign img[11544] = 77;
assign img[11545] = 81;
assign img[11546] = 80;
assign img[11547] = 79;
assign img[11548] = 76;
assign img[11549] = 81;
assign img[11550] = 79;
assign img[11551] = 77;
assign img[11552] = 81;
assign img[11553] = 75;
assign img[11554] = 81;
assign img[11555] = 72;
assign img[11556] = 77;
assign img[11557] = 75;
assign img[11558] = 76;
assign img[11559] = 77;
assign img[11560] = 72;
assign img[11561] = 73;
assign img[11562] = 82;
assign img[11563] = 84;
assign img[11564] = 84;
assign img[11565] = 73;
assign img[11566] = 78;
assign img[11567] = 76;
assign img[11568] = 80;
assign img[11569] = 76;
assign img[11570] = 80;
assign img[11571] = 84;
assign img[11572] = 80;
assign img[11573] = 74;
assign img[11574] = 81;
assign img[11575] = 77;
assign img[11576] = 77;
assign img[11577] = 77;
assign img[11578] = 81;
assign img[11579] = 78;
assign img[11580] = 80;
assign img[11581] = 71;
assign img[11582] = 82;
assign img[11583] = 80;
assign img[11584] = 73;
assign img[11585] = 76;
assign img[11586] = 73;
assign img[11587] = 81;
assign img[11588] = 77;
assign img[11589] = 80;
assign img[11590] = 85;
assign img[11591] = 79;
assign img[11592] = 70;
assign img[11593] = 75;
assign img[11594] = 73;
assign img[11595] = 69;
assign img[11596] = 72;
assign img[11597] = 73;
assign img[11598] = 72;
assign img[11599] = 66;
assign img[11600] = 65;
assign img[11601] = 64;
assign img[11602] = 64;
assign img[11603] = 59;
assign img[11604] = 56;
assign img[11605] = 49;
assign img[11606] = 53;
assign img[11607] = 56;
assign img[11608] = 51;
assign img[11609] = 54;
assign img[11610] = 56;
assign img[11611] = 56;
assign img[11612] = 50;
assign img[11613] = 52;
assign img[11614] = 53;
assign img[11615] = 49;
assign img[11616] = 48;
assign img[11617] = 54;
assign img[11618] = 50;
assign img[11619] = 51;
assign img[11620] = 47;
assign img[11621] = 53;
assign img[11622] = 48;
assign img[11623] = 56;
assign img[11624] = 50;
assign img[11625] = 49;
assign img[11626] = 50;
assign img[11627] = 52;
assign img[11628] = 51;
assign img[11629] = 53;
assign img[11630] = 48;
assign img[11631] = 47;
assign img[11632] = 49;
assign img[11633] = 51;
assign img[11634] = 48;
assign img[11635] = 52;
assign img[11636] = 56;
assign img[11637] = 50;
assign img[11638] = 48;
assign img[11639] = 48;
assign img[11640] = 46;
assign img[11641] = 45;
assign img[11642] = 44;
assign img[11643] = 49;
assign img[11644] = 50;
assign img[11645] = 49;
assign img[11646] = 49;
assign img[11647] = 48;
assign img[11648] = 48;
assign img[11649] = 42;
assign img[11650] = 45;
assign img[11651] = 47;
assign img[11652] = 46;
assign img[11653] = 52;
assign img[11654] = 55;
assign img[11655] = 64;
assign img[11656] = 68;
assign img[11657] = 65;
assign img[11658] = 64;
assign img[11659] = 65;
assign img[11660] = 64;
assign img[11661] = 64;
assign img[11662] = 64;
assign img[11663] = 65;
assign img[11664] = 69;
assign img[11665] = 68;
assign img[11666] = 66;
assign img[11667] = 66;
assign img[11668] = 66;
assign img[11669] = 69;
assign img[11670] = 64;
assign img[11671] = 65;
assign img[11672] = 65;
assign img[11673] = 64;
assign img[11674] = 66;
assign img[11675] = 69;
assign img[11676] = 65;
assign img[11677] = 65;
assign img[11678] = 65;
assign img[11679] = 73;
assign img[11680] = 64;
assign img[11681] = 69;
assign img[11682] = 65;
assign img[11683] = 67;
assign img[11684] = 65;
assign img[11685] = 65;
assign img[11686] = 66;
assign img[11687] = 65;
assign img[11688] = 67;
assign img[11689] = 65;
assign img[11690] = 70;
assign img[11691] = 76;
assign img[11692] = 70;
assign img[11693] = 64;
assign img[11694] = 67;
assign img[11695] = 73;
assign img[11696] = 64;
assign img[11697] = 68;
assign img[11698] = 64;
assign img[11699] = 65;
assign img[11700] = 65;
assign img[11701] = 72;
assign img[11702] = 64;
assign img[11703] = 65;
assign img[11704] = 64;
assign img[11705] = 66;
assign img[11706] = 64;
assign img[11707] = 70;
assign img[11708] = 65;
assign img[11709] = 66;
assign img[11710] = 70;
assign img[11711] = 65;
assign img[11712] = 64;
assign img[11713] = 67;
assign img[11714] = 64;
assign img[11715] = 65;
assign img[11716] = 67;
assign img[11717] = 64;
assign img[11718] = 68;
assign img[11719] = 66;
assign img[11720] = 68;
assign img[11721] = 64;
assign img[11722] = 64;
assign img[11723] = 64;
assign img[11724] = 64;
assign img[11725] = 64;
assign img[11726] = 64;
assign img[11727] = 53;
assign img[11728] = 51;
assign img[11729] = 42;
assign img[11730] = 49;
assign img[11731] = 44;
assign img[11732] = 46;
assign img[11733] = 45;
assign img[11734] = 44;
assign img[11735] = 41;
assign img[11736] = 38;
assign img[11737] = 43;
assign img[11738] = 41;
assign img[11739] = 39;
assign img[11740] = 38;
assign img[11741] = 44;
assign img[11742] = 39;
assign img[11743] = 36;
assign img[11744] = 39;
assign img[11745] = 39;
assign img[11746] = 44;
assign img[11747] = 37;
assign img[11748] = 42;
assign img[11749] = 41;
assign img[11750] = 36;
assign img[11751] = 41;
assign img[11752] = 41;
assign img[11753] = 39;
assign img[11754] = 37;
assign img[11755] = 49;
assign img[11756] = 33;
assign img[11757] = 38;
assign img[11758] = 40;
assign img[11759] = 45;
assign img[11760] = 44;
assign img[11761] = 35;
assign img[11762] = 37;
assign img[11763] = 33;
assign img[11764] = 36;
assign img[11765] = 38;
assign img[11766] = 38;
assign img[11767] = 36;
assign img[11768] = 36;
assign img[11769] = 38;
assign img[11770] = 33;
assign img[11771] = 34;
assign img[11772] = 37;
assign img[11773] = 38;
assign img[11774] = 40;
assign img[11775] = 40;
assign img[11776] = 44;
assign img[11777] = 50;
assign img[11778] = 52;
assign img[11779] = 51;
assign img[11780] = 54;
assign img[11781] = 48;
assign img[11782] = 64;
assign img[11783] = 66;
assign img[11784] = 69;
assign img[11785] = 72;
assign img[11786] = 65;
assign img[11787] = 64;
assign img[11788] = 68;
assign img[11789] = 64;
assign img[11790] = 65;
assign img[11791] = 65;
assign img[11792] = 66;
assign img[11793] = 68;
assign img[11794] = 65;
assign img[11795] = 70;
assign img[11796] = 65;
assign img[11797] = 65;
assign img[11798] = 66;
assign img[11799] = 64;
assign img[11800] = 67;
assign img[11801] = 64;
assign img[11802] = 65;
assign img[11803] = 65;
assign img[11804] = 65;
assign img[11805] = 66;
assign img[11806] = 73;
assign img[11807] = 69;
assign img[11808] = 72;
assign img[11809] = 67;
assign img[11810] = 68;
assign img[11811] = 68;
assign img[11812] = 66;
assign img[11813] = 69;
assign img[11814] = 68;
assign img[11815] = 67;
assign img[11816] = 64;
assign img[11817] = 69;
assign img[11818] = 65;
assign img[11819] = 68;
assign img[11820] = 77;
assign img[11821] = 69;
assign img[11822] = 72;
assign img[11823] = 65;
assign img[11824] = 70;
assign img[11825] = 68;
assign img[11826] = 68;
assign img[11827] = 65;
assign img[11828] = 65;
assign img[11829] = 65;
assign img[11830] = 71;
assign img[11831] = 76;
assign img[11832] = 69;
assign img[11833] = 65;
assign img[11834] = 65;
assign img[11835] = 68;
assign img[11836] = 73;
assign img[11837] = 65;
assign img[11838] = 64;
assign img[11839] = 70;
assign img[11840] = 65;
assign img[11841] = 65;
assign img[11842] = 70;
assign img[11843] = 78;
assign img[11844] = 66;
assign img[11845] = 67;
assign img[11846] = 67;
assign img[11847] = 72;
assign img[11848] = 68;
assign img[11849] = 70;
assign img[11850] = 69;
assign img[11851] = 65;
assign img[11852] = 68;
assign img[11853] = 66;
assign img[11854] = 65;
assign img[11855] = 64;
assign img[11856] = 52;
assign img[11857] = 48;
assign img[11858] = 48;
assign img[11859] = 50;
assign img[11860] = 52;
assign img[11861] = 46;
assign img[11862] = 48;
assign img[11863] = 52;
assign img[11864] = 44;
assign img[11865] = 48;
assign img[11866] = 45;
assign img[11867] = 46;
assign img[11868] = 44;
assign img[11869] = 46;
assign img[11870] = 46;
assign img[11871] = 45;
assign img[11872] = 39;
assign img[11873] = 47;
assign img[11874] = 41;
assign img[11875] = 48;
assign img[11876] = 38;
assign img[11877] = 42;
assign img[11878] = 44;
assign img[11879] = 44;
assign img[11880] = 42;
assign img[11881] = 36;
assign img[11882] = 44;
assign img[11883] = 44;
assign img[11884] = 44;
assign img[11885] = 40;
assign img[11886] = 46;
assign img[11887] = 39;
assign img[11888] = 38;
assign img[11889] = 42;
assign img[11890] = 39;
assign img[11891] = 46;
assign img[11892] = 38;
assign img[11893] = 40;
assign img[11894] = 44;
assign img[11895] = 39;
assign img[11896] = 38;
assign img[11897] = 44;
assign img[11898] = 44;
assign img[11899] = 42;
assign img[11900] = 39;
assign img[11901] = 49;
assign img[11902] = 46;
assign img[11903] = 44;
assign img[11904] = 44;
assign img[11905] = 43;
assign img[11906] = 44;
assign img[11907] = 44;
assign img[11908] = 41;
assign img[11909] = 54;
assign img[11910] = 50;
assign img[11911] = 56;
assign img[11912] = 64;
assign img[11913] = 65;
assign img[11914] = 64;
assign img[11915] = 64;
assign img[11916] = 64;
assign img[11917] = 69;
assign img[11918] = 64;
assign img[11919] = 64;
assign img[11920] = 64;
assign img[11921] = 65;
assign img[11922] = 68;
assign img[11923] = 65;
assign img[11924] = 64;
assign img[11925] = 66;
assign img[11926] = 67;
assign img[11927] = 65;
assign img[11928] = 64;
assign img[11929] = 65;
assign img[11930] = 65;
assign img[11931] = 65;
assign img[11932] = 67;
assign img[11933] = 64;
assign img[11934] = 64;
assign img[11935] = 67;
assign img[11936] = 72;
assign img[11937] = 69;
assign img[11938] = 72;
assign img[11939] = 65;
assign img[11940] = 65;
assign img[11941] = 64;
assign img[11942] = 69;
assign img[11943] = 70;
assign img[11944] = 65;
assign img[11945] = 65;
assign img[11946] = 66;
assign img[11947] = 64;
assign img[11948] = 65;
assign img[11949] = 67;
assign img[11950] = 65;
assign img[11951] = 67;
assign img[11952] = 67;
assign img[11953] = 64;
assign img[11954] = 64;
assign img[11955] = 70;
assign img[11956] = 70;
assign img[11957] = 69;
assign img[11958] = 65;
assign img[11959] = 57;
assign img[11960] = 67;
assign img[11961] = 64;
assign img[11962] = 67;
assign img[11963] = 65;
assign img[11964] = 66;
assign img[11965] = 69;
assign img[11966] = 65;
assign img[11967] = 73;
assign img[11968] = 65;
assign img[11969] = 66;
assign img[11970] = 65;
assign img[11971] = 65;
assign img[11972] = 66;
assign img[11973] = 73;
assign img[11974] = 66;
assign img[11975] = 68;
assign img[11976] = 64;
assign img[11977] = 65;
assign img[11978] = 65;
assign img[11979] = 64;
assign img[11980] = 65;
assign img[11981] = 64;
assign img[11982] = 64;
assign img[11983] = 64;
assign img[11984] = 56;
assign img[11985] = 42;
assign img[11986] = 40;
assign img[11987] = 46;
assign img[11988] = 50;
assign img[11989] = 44;
assign img[11990] = 46;
assign img[11991] = 44;
assign img[11992] = 37;
assign img[11993] = 40;
assign img[11994] = 39;
assign img[11995] = 41;
assign img[11996] = 39;
assign img[11997] = 40;
assign img[11998] = 36;
assign img[11999] = 42;
assign img[12000] = 36;
assign img[12001] = 37;
assign img[12002] = 38;
assign img[12003] = 37;
assign img[12004] = 38;
assign img[12005] = 39;
assign img[12006] = 36;
assign img[12007] = 41;
assign img[12008] = 40;
assign img[12009] = 35;
assign img[12010] = 32;
assign img[12011] = 33;
assign img[12012] = 34;
assign img[12013] = 36;
assign img[12014] = 33;
assign img[12015] = 41;
assign img[12016] = 39;
assign img[12017] = 34;
assign img[12018] = 35;
assign img[12019] = 37;
assign img[12020] = 35;
assign img[12021] = 32;
assign img[12022] = 28;
assign img[12023] = 34;
assign img[12024] = 43;
assign img[12025] = 38;
assign img[12026] = 32;
assign img[12027] = 36;
assign img[12028] = 38;
assign img[12029] = 37;
assign img[12030] = 33;
assign img[12031] = 36;
assign img[12032] = 36;
assign img[12033] = 64;
assign img[12034] = 64;
assign img[12035] = 64;
assign img[12036] = 64;
assign img[12037] = 65;
assign img[12038] = 66;
assign img[12039] = 68;
assign img[12040] = 73;
assign img[12041] = 78;
assign img[12042] = 73;
assign img[12043] = 81;
assign img[12044] = 73;
assign img[12045] = 69;
assign img[12046] = 73;
assign img[12047] = 78;
assign img[12048] = 73;
assign img[12049] = 69;
assign img[12050] = 75;
assign img[12051] = 73;
assign img[12052] = 70;
assign img[12053] = 75;
assign img[12054] = 68;
assign img[12055] = 74;
assign img[12056] = 81;
assign img[12057] = 73;
assign img[12058] = 72;
assign img[12059] = 76;
assign img[12060] = 74;
assign img[12061] = 71;
assign img[12062] = 77;
assign img[12063] = 73;
assign img[12064] = 72;
assign img[12065] = 73;
assign img[12066] = 73;
assign img[12067] = 74;
assign img[12068] = 74;
assign img[12069] = 72;
assign img[12070] = 69;
assign img[12071] = 71;
assign img[12072] = 78;
assign img[12073] = 77;
assign img[12074] = 78;
assign img[12075] = 73;
assign img[12076] = 77;
assign img[12077] = 73;
assign img[12078] = 78;
assign img[12079] = 84;
assign img[12080] = 76;
assign img[12081] = 68;
assign img[12082] = 69;
assign img[12083] = 77;
assign img[12084] = 73;
assign img[12085] = 77;
assign img[12086] = 76;
assign img[12087] = 73;
assign img[12088] = 72;
assign img[12089] = 70;
assign img[12090] = 77;
assign img[12091] = 78;
assign img[12092] = 77;
assign img[12093] = 72;
assign img[12094] = 73;
assign img[12095] = 77;
assign img[12096] = 77;
assign img[12097] = 77;
assign img[12098] = 73;
assign img[12099] = 77;
assign img[12100] = 80;
assign img[12101] = 77;
assign img[12102] = 77;
assign img[12103] = 73;
assign img[12104] = 77;
assign img[12105] = 73;
assign img[12106] = 69;
assign img[12107] = 70;
assign img[12108] = 74;
assign img[12109] = 73;
assign img[12110] = 78;
assign img[12111] = 72;
assign img[12112] = 65;
assign img[12113] = 64;
assign img[12114] = 52;
assign img[12115] = 64;
assign img[12116] = 53;
assign img[12117] = 52;
assign img[12118] = 52;
assign img[12119] = 64;
assign img[12120] = 48;
assign img[12121] = 60;
assign img[12122] = 52;
assign img[12123] = 56;
assign img[12124] = 54;
assign img[12125] = 54;
assign img[12126] = 44;
assign img[12127] = 46;
assign img[12128] = 52;
assign img[12129] = 52;
assign img[12130] = 51;
assign img[12131] = 47;
assign img[12132] = 46;
assign img[12133] = 44;
assign img[12134] = 44;
assign img[12135] = 46;
assign img[12136] = 45;
assign img[12137] = 46;
assign img[12138] = 46;
assign img[12139] = 41;
assign img[12140] = 42;
assign img[12141] = 44;
assign img[12142] = 42;
assign img[12143] = 45;
assign img[12144] = 44;
assign img[12145] = 44;
assign img[12146] = 44;
assign img[12147] = 44;
assign img[12148] = 44;
assign img[12149] = 44;
assign img[12150] = 47;
assign img[12151] = 44;
assign img[12152] = 45;
assign img[12153] = 46;
assign img[12154] = 44;
assign img[12155] = 44;
assign img[12156] = 44;
assign img[12157] = 42;
assign img[12158] = 47;
assign img[12159] = 44;
assign img[12160] = 45;
assign img[12161] = 46;
assign img[12162] = 48;
assign img[12163] = 52;
assign img[12164] = 48;
assign img[12165] = 49;
assign img[12166] = 49;
assign img[12167] = 64;
assign img[12168] = 65;
assign img[12169] = 67;
assign img[12170] = 65;
assign img[12171] = 65;
assign img[12172] = 64;
assign img[12173] = 69;
assign img[12174] = 65;
assign img[12175] = 64;
assign img[12176] = 66;
assign img[12177] = 69;
assign img[12178] = 57;
assign img[12179] = 67;
assign img[12180] = 73;
assign img[12181] = 64;
assign img[12182] = 64;
assign img[12183] = 66;
assign img[12184] = 67;
assign img[12185] = 65;
assign img[12186] = 69;
assign img[12187] = 68;
assign img[12188] = 64;
assign img[12189] = 66;
assign img[12190] = 64;
assign img[12191] = 65;
assign img[12192] = 65;
assign img[12193] = 65;
assign img[12194] = 64;
assign img[12195] = 64;
assign img[12196] = 66;
assign img[12197] = 65;
assign img[12198] = 64;
assign img[12199] = 66;
assign img[12200] = 65;
assign img[12201] = 65;
assign img[12202] = 64;
assign img[12203] = 57;
assign img[12204] = 68;
assign img[12205] = 65;
assign img[12206] = 64;
assign img[12207] = 73;
assign img[12208] = 65;
assign img[12209] = 64;
assign img[12210] = 64;
assign img[12211] = 66;
assign img[12212] = 65;
assign img[12213] = 64;
assign img[12214] = 66;
assign img[12215] = 64;
assign img[12216] = 64;
assign img[12217] = 65;
assign img[12218] = 69;
assign img[12219] = 64;
assign img[12220] = 65;
assign img[12221] = 64;
assign img[12222] = 65;
assign img[12223] = 64;
assign img[12224] = 65;
assign img[12225] = 69;
assign img[12226] = 64;
assign img[12227] = 67;
assign img[12228] = 66;
assign img[12229] = 64;
assign img[12230] = 64;
assign img[12231] = 65;
assign img[12232] = 55;
assign img[12233] = 64;
assign img[12234] = 69;
assign img[12235] = 57;
assign img[12236] = 65;
assign img[12237] = 64;
assign img[12238] = 70;
assign img[12239] = 65;
assign img[12240] = 67;
assign img[12241] = 57;
assign img[12242] = 51;
assign img[12243] = 48;
assign img[12244] = 42;
assign img[12245] = 42;
assign img[12246] = 50;
assign img[12247] = 42;
assign img[12248] = 41;
assign img[12249] = 43;
assign img[12250] = 40;
assign img[12251] = 46;
assign img[12252] = 43;
assign img[12253] = 45;
assign img[12254] = 45;
assign img[12255] = 38;
assign img[12256] = 45;
assign img[12257] = 41;
assign img[12258] = 41;
assign img[12259] = 41;
assign img[12260] = 37;
assign img[12261] = 42;
assign img[12262] = 36;
assign img[12263] = 39;
assign img[12264] = 41;
assign img[12265] = 40;
assign img[12266] = 34;
assign img[12267] = 44;
assign img[12268] = 41;
assign img[12269] = 40;
assign img[12270] = 42;
assign img[12271] = 38;
assign img[12272] = 34;
assign img[12273] = 40;
assign img[12274] = 40;
assign img[12275] = 37;
assign img[12276] = 37;
assign img[12277] = 33;
assign img[12278] = 39;
assign img[12279] = 41;
assign img[12280] = 37;
assign img[12281] = 37;
assign img[12282] = 35;
assign img[12283] = 38;
assign img[12284] = 40;
assign img[12285] = 37;
assign img[12286] = 36;
assign img[12287] = 38;
assign img[12288] = 64;
assign img[12289] = 40;
assign img[12290] = 37;
assign img[12291] = 40;
assign img[12292] = 39;
assign img[12293] = 47;
assign img[12294] = 46;
assign img[12295] = 46;
assign img[12296] = 48;
assign img[12297] = 55;
assign img[12298] = 64;
assign img[12299] = 65;
assign img[12300] = 53;
assign img[12301] = 64;
assign img[12302] = 55;
assign img[12303] = 55;
assign img[12304] = 64;
assign img[12305] = 54;
assign img[12306] = 55;
assign img[12307] = 56;
assign img[12308] = 64;
assign img[12309] = 64;
assign img[12310] = 64;
assign img[12311] = 53;
assign img[12312] = 64;
assign img[12313] = 54;
assign img[12314] = 64;
assign img[12315] = 64;
assign img[12316] = 54;
assign img[12317] = 50;
assign img[12318] = 56;
assign img[12319] = 64;
assign img[12320] = 64;
assign img[12321] = 57;
assign img[12322] = 66;
assign img[12323] = 64;
assign img[12324] = 55;
assign img[12325] = 55;
assign img[12326] = 64;
assign img[12327] = 64;
assign img[12328] = 64;
assign img[12329] = 52;
assign img[12330] = 54;
assign img[12331] = 64;
assign img[12332] = 64;
assign img[12333] = 57;
assign img[12334] = 56;
assign img[12335] = 59;
assign img[12336] = 60;
assign img[12337] = 64;
assign img[12338] = 55;
assign img[12339] = 64;
assign img[12340] = 64;
assign img[12341] = 64;
assign img[12342] = 57;
assign img[12343] = 58;
assign img[12344] = 54;
assign img[12345] = 64;
assign img[12346] = 58;
assign img[12347] = 64;
assign img[12348] = 56;
assign img[12349] = 55;
assign img[12350] = 66;
assign img[12351] = 64;
assign img[12352] = 56;
assign img[12353] = 58;
assign img[12354] = 58;
assign img[12355] = 66;
assign img[12356] = 64;
assign img[12357] = 54;
assign img[12358] = 59;
assign img[12359] = 64;
assign img[12360] = 64;
assign img[12361] = 64;
assign img[12362] = 55;
assign img[12363] = 64;
assign img[12364] = 58;
assign img[12365] = 56;
assign img[12366] = 53;
assign img[12367] = 64;
assign img[12368] = 54;
assign img[12369] = 50;
assign img[12370] = 46;
assign img[12371] = 48;
assign img[12372] = 44;
assign img[12373] = 41;
assign img[12374] = 38;
assign img[12375] = 44;
assign img[12376] = 44;
assign img[12377] = 36;
assign img[12378] = 39;
assign img[12379] = 39;
assign img[12380] = 38;
assign img[12381] = 36;
assign img[12382] = 36;
assign img[12383] = 37;
assign img[12384] = 33;
assign img[12385] = 38;
assign img[12386] = 32;
assign img[12387] = 36;
assign img[12388] = 36;
assign img[12389] = 36;
assign img[12390] = 33;
assign img[12391] = 29;
assign img[12392] = 34;
assign img[12393] = 36;
assign img[12394] = 32;
assign img[12395] = 32;
assign img[12396] = 32;
assign img[12397] = 36;
assign img[12398] = 34;
assign img[12399] = 34;
assign img[12400] = 30;
assign img[12401] = 32;
assign img[12402] = 32;
assign img[12403] = 32;
assign img[12404] = 32;
assign img[12405] = 32;
assign img[12406] = 32;
assign img[12407] = 32;
assign img[12408] = 28;
assign img[12409] = 34;
assign img[12410] = 28;
assign img[12411] = 34;
assign img[12412] = 32;
assign img[12413] = 32;
assign img[12414] = 28;
assign img[12415] = 34;
assign img[12416] = 28;
assign img[12417] = 70;
assign img[12418] = 74;
assign img[12419] = 68;
assign img[12420] = 68;
assign img[12421] = 72;
assign img[12422] = 74;
assign img[12423] = 76;
assign img[12424] = 77;
assign img[12425] = 76;
assign img[12426] = 78;
assign img[12427] = 85;
assign img[12428] = 86;
assign img[12429] = 87;
assign img[12430] = 86;
assign img[12431] = 81;
assign img[12432] = 90;
assign img[12433] = 94;
assign img[12434] = 88;
assign img[12435] = 88;
assign img[12436] = 88;
assign img[12437] = 88;
assign img[12438] = 92;
assign img[12439] = 87;
assign img[12440] = 88;
assign img[12441] = 88;
assign img[12442] = 87;
assign img[12443] = 80;
assign img[12444] = 87;
assign img[12445] = 88;
assign img[12446] = 87;
assign img[12447] = 88;
assign img[12448] = 87;
assign img[12449] = 94;
assign img[12450] = 96;
assign img[12451] = 92;
assign img[12452] = 84;
assign img[12453] = 85;
assign img[12454] = 88;
assign img[12455] = 88;
assign img[12456] = 86;
assign img[12457] = 94;
assign img[12458] = 88;
assign img[12459] = 80;
assign img[12460] = 88;
assign img[12461] = 87;
assign img[12462] = 94;
assign img[12463] = 87;
assign img[12464] = 87;
assign img[12465] = 94;
assign img[12466] = 87;
assign img[12467] = 98;
assign img[12468] = 87;
assign img[12469] = 88;
assign img[12470] = 94;
assign img[12471] = 88;
assign img[12472] = 88;
assign img[12473] = 92;
assign img[12474] = 84;
assign img[12475] = 86;
assign img[12476] = 84;
assign img[12477] = 84;
assign img[12478] = 77;
assign img[12479] = 81;
assign img[12480] = 84;
assign img[12481] = 85;
assign img[12482] = 84;
assign img[12483] = 86;
assign img[12484] = 76;
assign img[12485] = 80;
assign img[12486] = 82;
assign img[12487] = 84;
assign img[12488] = 81;
assign img[12489] = 84;
assign img[12490] = 84;
assign img[12491] = 85;
assign img[12492] = 79;
assign img[12493] = 78;
assign img[12494] = 86;
assign img[12495] = 79;
assign img[12496] = 84;
assign img[12497] = 83;
assign img[12498] = 80;
assign img[12499] = 78;
assign img[12500] = 78;
assign img[12501] = 70;
assign img[12502] = 66;
assign img[12503] = 70;
assign img[12504] = 64;
assign img[12505] = 64;
assign img[12506] = 72;
assign img[12507] = 68;
assign img[12508] = 64;
assign img[12509] = 64;
assign img[12510] = 68;
assign img[12511] = 65;
assign img[12512] = 64;
assign img[12513] = 64;
assign img[12514] = 64;
assign img[12515] = 64;
assign img[12516] = 60;
assign img[12517] = 64;
assign img[12518] = 64;
assign img[12519] = 64;
assign img[12520] = 56;
assign img[12521] = 56;
assign img[12522] = 68;
assign img[12523] = 58;
assign img[12524] = 64;
assign img[12525] = 64;
assign img[12526] = 60;
assign img[12527] = 55;
assign img[12528] = 64;
assign img[12529] = 64;
assign img[12530] = 64;
assign img[12531] = 56;
assign img[12532] = 60;
assign img[12533] = 53;
assign img[12534] = 64;
assign img[12535] = 52;
assign img[12536] = 56;
assign img[12537] = 60;
assign img[12538] = 52;
assign img[12539] = 56;
assign img[12540] = 55;
assign img[12541] = 59;
assign img[12542] = 64;
assign img[12543] = 64;
assign img[12544] = 64;
assign img[12545] = 32;
assign img[12546] = 36;
assign img[12547] = 32;
assign img[12548] = 44;
assign img[12549] = 36;
assign img[12550] = 40;
assign img[12551] = 46;
assign img[12552] = 45;
assign img[12553] = 52;
assign img[12554] = 50;
assign img[12555] = 53;
assign img[12556] = 55;
assign img[12557] = 48;
assign img[12558] = 52;
assign img[12559] = 55;
assign img[12560] = 64;
assign img[12561] = 55;
assign img[12562] = 55;
assign img[12563] = 54;
assign img[12564] = 53;
assign img[12565] = 53;
assign img[12566] = 48;
assign img[12567] = 55;
assign img[12568] = 48;
assign img[12569] = 54;
assign img[12570] = 51;
assign img[12571] = 55;
assign img[12572] = 56;
assign img[12573] = 54;
assign img[12574] = 56;
assign img[12575] = 60;
assign img[12576] = 53;
assign img[12577] = 56;
assign img[12578] = 57;
assign img[12579] = 54;
assign img[12580] = 46;
assign img[12581] = 49;
assign img[12582] = 64;
assign img[12583] = 64;
assign img[12584] = 60;
assign img[12585] = 54;
assign img[12586] = 48;
assign img[12587] = 64;
assign img[12588] = 55;
assign img[12589] = 51;
assign img[12590] = 44;
assign img[12591] = 58;
assign img[12592] = 52;
assign img[12593] = 47;
assign img[12594] = 54;
assign img[12595] = 48;
assign img[12596] = 54;
assign img[12597] = 55;
assign img[12598] = 56;
assign img[12599] = 53;
assign img[12600] = 56;
assign img[12601] = 60;
assign img[12602] = 54;
assign img[12603] = 57;
assign img[12604] = 51;
assign img[12605] = 64;
assign img[12606] = 55;
assign img[12607] = 48;
assign img[12608] = 53;
assign img[12609] = 53;
assign img[12610] = 53;
assign img[12611] = 51;
assign img[12612] = 47;
assign img[12613] = 52;
assign img[12614] = 53;
assign img[12615] = 53;
assign img[12616] = 49;
assign img[12617] = 52;
assign img[12618] = 53;
assign img[12619] = 51;
assign img[12620] = 56;
assign img[12621] = 56;
assign img[12622] = 56;
assign img[12623] = 52;
assign img[12624] = 48;
assign img[12625] = 50;
assign img[12626] = 48;
assign img[12627] = 48;
assign img[12628] = 43;
assign img[12629] = 44;
assign img[12630] = 41;
assign img[12631] = 36;
assign img[12632] = 28;
assign img[12633] = 35;
assign img[12634] = 30;
assign img[12635] = 36;
assign img[12636] = 30;
assign img[12637] = 29;
assign img[12638] = 30;
assign img[12639] = 24;
assign img[12640] = 34;
assign img[12641] = 32;
assign img[12642] = 34;
assign img[12643] = 30;
assign img[12644] = 28;
assign img[12645] = 27;
assign img[12646] = 25;
assign img[12647] = 30;
assign img[12648] = 32;
assign img[12649] = 29;
assign img[12650] = 30;
assign img[12651] = 25;
assign img[12652] = 29;
assign img[12653] = 25;
assign img[12654] = 29;
assign img[12655] = 28;
assign img[12656] = 23;
assign img[12657] = 26;
assign img[12658] = 25;
assign img[12659] = 25;
assign img[12660] = 31;
assign img[12661] = 22;
assign img[12662] = 28;
assign img[12663] = 24;
assign img[12664] = 28;
assign img[12665] = 25;
assign img[12666] = 27;
assign img[12667] = 25;
assign img[12668] = 26;
assign img[12669] = 21;
assign img[12670] = 24;
assign img[12671] = 23;
assign img[12672] = 27;
assign img[12673] = 34;
assign img[12674] = 34;
assign img[12675] = 34;
assign img[12676] = 33;
assign img[12677] = 29;
assign img[12678] = 34;
assign img[12679] = 40;
assign img[12680] = 42;
assign img[12681] = 42;
assign img[12682] = 42;
assign img[12683] = 47;
assign img[12684] = 46;
assign img[12685] = 50;
assign img[12686] = 48;
assign img[12687] = 48;
assign img[12688] = 52;
assign img[12689] = 46;
assign img[12690] = 50;
assign img[12691] = 49;
assign img[12692] = 48;
assign img[12693] = 46;
assign img[12694] = 48;
assign img[12695] = 52;
assign img[12696] = 44;
assign img[12697] = 48;
assign img[12698] = 54;
assign img[12699] = 54;
assign img[12700] = 40;
assign img[12701] = 51;
assign img[12702] = 50;
assign img[12703] = 52;
assign img[12704] = 47;
assign img[12705] = 48;
assign img[12706] = 50;
assign img[12707] = 48;
assign img[12708] = 46;
assign img[12709] = 48;
assign img[12710] = 47;
assign img[12711] = 48;
assign img[12712] = 54;
assign img[12713] = 52;
assign img[12714] = 50;
assign img[12715] = 64;
assign img[12716] = 48;
assign img[12717] = 47;
assign img[12718] = 46;
assign img[12719] = 54;
assign img[12720] = 50;
assign img[12721] = 47;
assign img[12722] = 50;
assign img[12723] = 44;
assign img[12724] = 46;
assign img[12725] = 46;
assign img[12726] = 39;
assign img[12727] = 47;
assign img[12728] = 44;
assign img[12729] = 54;
assign img[12730] = 54;
assign img[12731] = 48;
assign img[12732] = 46;
assign img[12733] = 48;
assign img[12734] = 51;
assign img[12735] = 50;
assign img[12736] = 41;
assign img[12737] = 40;
assign img[12738] = 44;
assign img[12739] = 48;
assign img[12740] = 53;
assign img[12741] = 45;
assign img[12742] = 50;
assign img[12743] = 45;
assign img[12744] = 40;
assign img[12745] = 45;
assign img[12746] = 56;
assign img[12747] = 49;
assign img[12748] = 42;
assign img[12749] = 57;
assign img[12750] = 42;
assign img[12751] = 48;
assign img[12752] = 43;
assign img[12753] = 50;
assign img[12754] = 49;
assign img[12755] = 48;
assign img[12756] = 41;
assign img[12757] = 37;
assign img[12758] = 38;
assign img[12759] = 34;
assign img[12760] = 26;
assign img[12761] = 28;
assign img[12762] = 28;
assign img[12763] = 28;
assign img[12764] = 33;
assign img[12765] = 32;
assign img[12766] = 30;
assign img[12767] = 26;
assign img[12768] = 30;
assign img[12769] = 32;
assign img[12770] = 26;
assign img[12771] = 27;
assign img[12772] = 29;
assign img[12773] = 25;
assign img[12774] = 26;
assign img[12775] = 27;
assign img[12776] = 26;
assign img[12777] = 28;
assign img[12778] = 24;
assign img[12779] = 25;
assign img[12780] = 24;
assign img[12781] = 19;
assign img[12782] = 25;
assign img[12783] = 27;
assign img[12784] = 24;
assign img[12785] = 25;
assign img[12786] = 22;
assign img[12787] = 28;
assign img[12788] = 20;
assign img[12789] = 21;
assign img[12790] = 19;
assign img[12791] = 19;
assign img[12792] = 22;
assign img[12793] = 20;
assign img[12794] = 24;
assign img[12795] = 24;
assign img[12796] = 21;
assign img[12797] = 18;
assign img[12798] = 22;
assign img[12799] = 26;
assign img[12800] = 18;
assign img[12801] = 55;
assign img[12802] = 56;
assign img[12803] = 57;
assign img[12804] = 50;
assign img[12805] = 57;
assign img[12806] = 64;
assign img[12807] = 64;
assign img[12808] = 65;
assign img[12809] = 68;
assign img[12810] = 64;
assign img[12811] = 73;
assign img[12812] = 70;
assign img[12813] = 71;
assign img[12814] = 68;
assign img[12815] = 68;
assign img[12816] = 76;
assign img[12817] = 78;
assign img[12818] = 71;
assign img[12819] = 79;
assign img[12820] = 76;
assign img[12821] = 72;
assign img[12822] = 72;
assign img[12823] = 72;
assign img[12824] = 70;
assign img[12825] = 76;
assign img[12826] = 78;
assign img[12827] = 65;
assign img[12828] = 77;
assign img[12829] = 70;
assign img[12830] = 70;
assign img[12831] = 76;
assign img[12832] = 73;
assign img[12833] = 72;
assign img[12834] = 70;
assign img[12835] = 77;
assign img[12836] = 72;
assign img[12837] = 80;
assign img[12838] = 70;
assign img[12839] = 76;
assign img[12840] = 72;
assign img[12841] = 78;
assign img[12842] = 71;
assign img[12843] = 74;
assign img[12844] = 71;
assign img[12845] = 70;
assign img[12846] = 69;
assign img[12847] = 69;
assign img[12848] = 72;
assign img[12849] = 70;
assign img[12850] = 78;
assign img[12851] = 71;
assign img[12852] = 70;
assign img[12853] = 74;
assign img[12854] = 72;
assign img[12855] = 69;
assign img[12856] = 70;
assign img[12857] = 76;
assign img[12858] = 68;
assign img[12859] = 71;
assign img[12860] = 64;
assign img[12861] = 65;
assign img[12862] = 68;
assign img[12863] = 69;
assign img[12864] = 69;
assign img[12865] = 72;
assign img[12866] = 72;
assign img[12867] = 72;
assign img[12868] = 68;
assign img[12869] = 68;
assign img[12870] = 68;
assign img[12871] = 65;
assign img[12872] = 70;
assign img[12873] = 68;
assign img[12874] = 65;
assign img[12875] = 73;
assign img[12876] = 68;
assign img[12877] = 65;
assign img[12878] = 69;
assign img[12879] = 66;
assign img[12880] = 66;
assign img[12881] = 66;
assign img[12882] = 69;
assign img[12883] = 67;
assign img[12884] = 66;
assign img[12885] = 66;
assign img[12886] = 64;
assign img[12887] = 51;
assign img[12888] = 52;
assign img[12889] = 52;
assign img[12890] = 53;
assign img[12891] = 50;
assign img[12892] = 57;
assign img[12893] = 48;
assign img[12894] = 50;
assign img[12895] = 58;
assign img[12896] = 49;
assign img[12897] = 49;
assign img[12898] = 48;
assign img[12899] = 51;
assign img[12900] = 53;
assign img[12901] = 49;
assign img[12902] = 47;
assign img[12903] = 45;
assign img[12904] = 49;
assign img[12905] = 46;
assign img[12906] = 47;
assign img[12907] = 46;
assign img[12908] = 46;
assign img[12909] = 44;
assign img[12910] = 48;
assign img[12911] = 41;
assign img[12912] = 47;
assign img[12913] = 43;
assign img[12914] = 40;
assign img[12915] = 41;
assign img[12916] = 41;
assign img[12917] = 45;
assign img[12918] = 43;
assign img[12919] = 36;
assign img[12920] = 44;
assign img[12921] = 43;
assign img[12922] = 46;
assign img[12923] = 46;
assign img[12924] = 40;
assign img[12925] = 45;
assign img[12926] = 44;
assign img[12927] = 46;
assign img[12928] = 42;
assign img[12929] = 40;
assign img[12930] = 33;
assign img[12931] = 38;
assign img[12932] = 40;
assign img[12933] = 40;
assign img[12934] = 49;
assign img[12935] = 44;
assign img[12936] = 44;
assign img[12937] = 52;
assign img[12938] = 50;
assign img[12939] = 54;
assign img[12940] = 64;
assign img[12941] = 55;
assign img[12942] = 52;
assign img[12943] = 64;
assign img[12944] = 52;
assign img[12945] = 55;
assign img[12946] = 54;
assign img[12947] = 55;
assign img[12948] = 64;
assign img[12949] = 53;
assign img[12950] = 64;
assign img[12951] = 54;
assign img[12952] = 52;
assign img[12953] = 47;
assign img[12954] = 55;
assign img[12955] = 64;
assign img[12956] = 52;
assign img[12957] = 56;
assign img[12958] = 55;
assign img[12959] = 54;
assign img[12960] = 64;
assign img[12961] = 55;
assign img[12962] = 56;
assign img[12963] = 54;
assign img[12964] = 54;
assign img[12965] = 56;
assign img[12966] = 55;
assign img[12967] = 54;
assign img[12968] = 56;
assign img[12969] = 55;
assign img[12970] = 64;
assign img[12971] = 52;
assign img[12972] = 51;
assign img[12973] = 56;
assign img[12974] = 54;
assign img[12975] = 64;
assign img[12976] = 55;
assign img[12977] = 53;
assign img[12978] = 55;
assign img[12979] = 64;
assign img[12980] = 54;
assign img[12981] = 55;
assign img[12982] = 54;
assign img[12983] = 51;
assign img[12984] = 64;
assign img[12985] = 64;
assign img[12986] = 54;
assign img[12987] = 64;
assign img[12988] = 64;
assign img[12989] = 55;
assign img[12990] = 50;
assign img[12991] = 48;
assign img[12992] = 50;
assign img[12993] = 51;
assign img[12994] = 51;
assign img[12995] = 56;
assign img[12996] = 53;
assign img[12997] = 51;
assign img[12998] = 48;
assign img[12999] = 50;
assign img[13000] = 52;
assign img[13001] = 52;
assign img[13002] = 52;
assign img[13003] = 50;
assign img[13004] = 48;
assign img[13005] = 52;
assign img[13006] = 47;
assign img[13007] = 52;
assign img[13008] = 46;
assign img[13009] = 50;
assign img[13010] = 46;
assign img[13011] = 45;
assign img[13012] = 50;
assign img[13013] = 52;
assign img[13014] = 41;
assign img[13015] = 40;
assign img[13016] = 36;
assign img[13017] = 33;
assign img[13018] = 38;
assign img[13019] = 35;
assign img[13020] = 36;
assign img[13021] = 33;
assign img[13022] = 36;
assign img[13023] = 35;
assign img[13024] = 36;
assign img[13025] = 32;
assign img[13026] = 29;
assign img[13027] = 37;
assign img[13028] = 34;
assign img[13029] = 33;
assign img[13030] = 34;
assign img[13031] = 32;
assign img[13032] = 34;
assign img[13033] = 33;
assign img[13034] = 33;
assign img[13035] = 29;
assign img[13036] = 30;
assign img[13037] = 30;
assign img[13038] = 32;
assign img[13039] = 32;
assign img[13040] = 32;
assign img[13041] = 30;
assign img[13042] = 26;
assign img[13043] = 32;
assign img[13044] = 29;
assign img[13045] = 32;
assign img[13046] = 28;
assign img[13047] = 28;
assign img[13048] = 31;
assign img[13049] = 30;
assign img[13050] = 32;
assign img[13051] = 28;
assign img[13052] = 32;
assign img[13053] = 32;
assign img[13054] = 27;
assign img[13055] = 30;
assign img[13056] = 28;
assign img[13057] = 37;
assign img[13058] = 33;
assign img[13059] = 35;
assign img[13060] = 38;
assign img[13061] = 40;
assign img[13062] = 42;
assign img[13063] = 38;
assign img[13064] = 47;
assign img[13065] = 41;
assign img[13066] = 52;
assign img[13067] = 54;
assign img[13068] = 52;
assign img[13069] = 51;
assign img[13070] = 64;
assign img[13071] = 50;
assign img[13072] = 57;
assign img[13073] = 52;
assign img[13074] = 46;
assign img[13075] = 50;
assign img[13076] = 52;
assign img[13077] = 56;
assign img[13078] = 50;
assign img[13079] = 50;
assign img[13080] = 49;
assign img[13081] = 49;
assign img[13082] = 55;
assign img[13083] = 56;
assign img[13084] = 52;
assign img[13085] = 53;
assign img[13086] = 53;
assign img[13087] = 52;
assign img[13088] = 52;
assign img[13089] = 51;
assign img[13090] = 57;
assign img[13091] = 54;
assign img[13092] = 57;
assign img[13093] = 56;
assign img[13094] = 50;
assign img[13095] = 64;
assign img[13096] = 53;
assign img[13097] = 49;
assign img[13098] = 57;
assign img[13099] = 56;
assign img[13100] = 56;
assign img[13101] = 52;
assign img[13102] = 53;
assign img[13103] = 48;
assign img[13104] = 54;
assign img[13105] = 46;
assign img[13106] = 52;
assign img[13107] = 53;
assign img[13108] = 50;
assign img[13109] = 53;
assign img[13110] = 49;
assign img[13111] = 53;
assign img[13112] = 53;
assign img[13113] = 52;
assign img[13114] = 49;
assign img[13115] = 54;
assign img[13116] = 56;
assign img[13117] = 51;
assign img[13118] = 51;
assign img[13119] = 50;
assign img[13120] = 53;
assign img[13121] = 52;
assign img[13122] = 54;
assign img[13123] = 53;
assign img[13124] = 55;
assign img[13125] = 54;
assign img[13126] = 53;
assign img[13127] = 52;
assign img[13128] = 49;
assign img[13129] = 54;
assign img[13130] = 49;
assign img[13131] = 50;
assign img[13132] = 56;
assign img[13133] = 49;
assign img[13134] = 52;
assign img[13135] = 48;
assign img[13136] = 51;
assign img[13137] = 50;
assign img[13138] = 47;
assign img[13139] = 46;
assign img[13140] = 50;
assign img[13141] = 44;
assign img[13142] = 49;
assign img[13143] = 45;
assign img[13144] = 38;
assign img[13145] = 39;
assign img[13146] = 36;
assign img[13147] = 34;
assign img[13148] = 32;
assign img[13149] = 39;
assign img[13150] = 32;
assign img[13151] = 33;
assign img[13152] = 33;
assign img[13153] = 33;
assign img[13154] = 33;
assign img[13155] = 36;
assign img[13156] = 30;
assign img[13157] = 34;
assign img[13158] = 36;
assign img[13159] = 32;
assign img[13160] = 32;
assign img[13161] = 29;
assign img[13162] = 28;
assign img[13163] = 32;
assign img[13164] = 34;
assign img[13165] = 33;
assign img[13166] = 32;
assign img[13167] = 29;
assign img[13168] = 32;
assign img[13169] = 26;
assign img[13170] = 30;
assign img[13171] = 34;
assign img[13172] = 25;
assign img[13173] = 25;
assign img[13174] = 26;
assign img[13175] = 32;
assign img[13176] = 29;
assign img[13177] = 32;
assign img[13178] = 32;
assign img[13179] = 25;
assign img[13180] = 26;
assign img[13181] = 29;
assign img[13182] = 34;
assign img[13183] = 26;
assign img[13184] = 30;
assign img[13185] = 56;
assign img[13186] = 53;
assign img[13187] = 47;
assign img[13188] = 58;
assign img[13189] = 64;
assign img[13190] = 64;
assign img[13191] = 57;
assign img[13192] = 64;
assign img[13193] = 64;
assign img[13194] = 68;
assign img[13195] = 66;
assign img[13196] = 65;
assign img[13197] = 65;
assign img[13198] = 65;
assign img[13199] = 73;
assign img[13200] = 73;
assign img[13201] = 69;
assign img[13202] = 73;
assign img[13203] = 68;
assign img[13204] = 68;
assign img[13205] = 70;
assign img[13206] = 67;
assign img[13207] = 69;
assign img[13208] = 69;
assign img[13209] = 69;
assign img[13210] = 73;
assign img[13211] = 71;
assign img[13212] = 70;
assign img[13213] = 73;
assign img[13214] = 69;
assign img[13215] = 68;
assign img[13216] = 69;
assign img[13217] = 73;
assign img[13218] = 65;
assign img[13219] = 69;
assign img[13220] = 69;
assign img[13221] = 68;
assign img[13222] = 69;
assign img[13223] = 69;
assign img[13224] = 66;
assign img[13225] = 68;
assign img[13226] = 70;
assign img[13227] = 67;
assign img[13228] = 65;
assign img[13229] = 68;
assign img[13230] = 69;
assign img[13231] = 73;
assign img[13232] = 65;
assign img[13233] = 73;
assign img[13234] = 69;
assign img[13235] = 65;
assign img[13236] = 64;
assign img[13237] = 65;
assign img[13238] = 65;
assign img[13239] = 66;
assign img[13240] = 67;
assign img[13241] = 77;
assign img[13242] = 76;
assign img[13243] = 73;
assign img[13244] = 67;
assign img[13245] = 69;
assign img[13246] = 73;
assign img[13247] = 69;
assign img[13248] = 69;
assign img[13249] = 71;
assign img[13250] = 64;
assign img[13251] = 65;
assign img[13252] = 73;
assign img[13253] = 69;
assign img[13254] = 73;
assign img[13255] = 73;
assign img[13256] = 65;
assign img[13257] = 64;
assign img[13258] = 73;
assign img[13259] = 65;
assign img[13260] = 65;
assign img[13261] = 65;
assign img[13262] = 65;
assign img[13263] = 65;
assign img[13264] = 65;
assign img[13265] = 72;
assign img[13266] = 64;
assign img[13267] = 66;
assign img[13268] = 64;
assign img[13269] = 65;
assign img[13270] = 65;
assign img[13271] = 64;
assign img[13272] = 64;
assign img[13273] = 49;
assign img[13274] = 52;
assign img[13275] = 47;
assign img[13276] = 47;
assign img[13277] = 52;
assign img[13278] = 48;
assign img[13279] = 49;
assign img[13280] = 48;
assign img[13281] = 52;
assign img[13282] = 45;
assign img[13283] = 46;
assign img[13284] = 44;
assign img[13285] = 47;
assign img[13286] = 44;
assign img[13287] = 43;
assign img[13288] = 47;
assign img[13289] = 47;
assign img[13290] = 48;
assign img[13291] = 45;
assign img[13292] = 47;
assign img[13293] = 41;
assign img[13294] = 47;
assign img[13295] = 45;
assign img[13296] = 48;
assign img[13297] = 44;
assign img[13298] = 45;
assign img[13299] = 44;
assign img[13300] = 45;
assign img[13301] = 44;
assign img[13302] = 44;
assign img[13303] = 44;
assign img[13304] = 41;
assign img[13305] = 45;
assign img[13306] = 41;
assign img[13307] = 48;
assign img[13308] = 47;
assign img[13309] = 44;
assign img[13310] = 44;
assign img[13311] = 37;
assign img[13312] = 41;
assign img[13313] = 46;
assign img[13314] = 38;
assign img[13315] = 43;
assign img[13316] = 44;
assign img[13317] = 44;
assign img[13318] = 48;
assign img[13319] = 45;
assign img[13320] = 52;
assign img[13321] = 53;
assign img[13322] = 50;
assign img[13323] = 64;
assign img[13324] = 54;
assign img[13325] = 56;
assign img[13326] = 64;
assign img[13327] = 64;
assign img[13328] = 57;
assign img[13329] = 53;
assign img[13330] = 64;
assign img[13331] = 64;
assign img[13332] = 56;
assign img[13333] = 64;
assign img[13334] = 64;
assign img[13335] = 57;
assign img[13336] = 58;
assign img[13337] = 54;
assign img[13338] = 64;
assign img[13339] = 64;
assign img[13340] = 55;
assign img[13341] = 64;
assign img[13342] = 53;
assign img[13343] = 65;
assign img[13344] = 64;
assign img[13345] = 64;
assign img[13346] = 57;
assign img[13347] = 56;
assign img[13348] = 64;
assign img[13349] = 53;
assign img[13350] = 64;
assign img[13351] = 64;
assign img[13352] = 53;
assign img[13353] = 56;
assign img[13354] = 64;
assign img[13355] = 64;
assign img[13356] = 53;
assign img[13357] = 56;
assign img[13358] = 56;
assign img[13359] = 58;
assign img[13360] = 64;
assign img[13361] = 55;
assign img[13362] = 64;
assign img[13363] = 51;
assign img[13364] = 64;
assign img[13365] = 64;
assign img[13366] = 53;
assign img[13367] = 52;
assign img[13368] = 64;
assign img[13369] = 64;
assign img[13370] = 57;
assign img[13371] = 64;
assign img[13372] = 64;
assign img[13373] = 56;
assign img[13374] = 56;
assign img[13375] = 56;
assign img[13376] = 64;
assign img[13377] = 64;
assign img[13378] = 57;
assign img[13379] = 64;
assign img[13380] = 57;
assign img[13381] = 58;
assign img[13382] = 58;
assign img[13383] = 52;
assign img[13384] = 52;
assign img[13385] = 64;
assign img[13386] = 64;
assign img[13387] = 56;
assign img[13388] = 56;
assign img[13389] = 64;
assign img[13390] = 64;
assign img[13391] = 55;
assign img[13392] = 64;
assign img[13393] = 54;
assign img[13394] = 52;
assign img[13395] = 55;
assign img[13396] = 51;
assign img[13397] = 56;
assign img[13398] = 51;
assign img[13399] = 54;
assign img[13400] = 48;
assign img[13401] = 46;
assign img[13402] = 42;
assign img[13403] = 38;
assign img[13404] = 39;
assign img[13405] = 40;
assign img[13406] = 39;
assign img[13407] = 40;
assign img[13408] = 38;
assign img[13409] = 36;
assign img[13410] = 44;
assign img[13411] = 39;
assign img[13412] = 40;
assign img[13413] = 39;
assign img[13414] = 38;
assign img[13415] = 37;
assign img[13416] = 41;
assign img[13417] = 41;
assign img[13418] = 39;
assign img[13419] = 37;
assign img[13420] = 36;
assign img[13421] = 38;
assign img[13422] = 34;
assign img[13423] = 38;
assign img[13424] = 33;
assign img[13425] = 34;
assign img[13426] = 37;
assign img[13427] = 39;
assign img[13428] = 33;
assign img[13429] = 33;
assign img[13430] = 36;
assign img[13431] = 35;
assign img[13432] = 33;
assign img[13433] = 32;
assign img[13434] = 34;
assign img[13435] = 37;
assign img[13436] = 34;
assign img[13437] = 32;
assign img[13438] = 29;
assign img[13439] = 32;
assign img[13440] = 32;
assign img[13441] = 52;
assign img[13442] = 50;
assign img[13443] = 49;
assign img[13444] = 50;
assign img[13445] = 48;
assign img[13446] = 64;
assign img[13447] = 64;
assign img[13448] = 64;
assign img[13449] = 64;
assign img[13450] = 64;
assign img[13451] = 65;
assign img[13452] = 64;
assign img[13453] = 68;
assign img[13454] = 56;
assign img[13455] = 64;
assign img[13456] = 64;
assign img[13457] = 65;
assign img[13458] = 68;
assign img[13459] = 64;
assign img[13460] = 64;
assign img[13461] = 68;
assign img[13462] = 69;
assign img[13463] = 64;
assign img[13464] = 64;
assign img[13465] = 65;
assign img[13466] = 68;
assign img[13467] = 70;
assign img[13468] = 64;
assign img[13469] = 64;
assign img[13470] = 68;
assign img[13471] = 64;
assign img[13472] = 64;
assign img[13473] = 64;
assign img[13474] = 73;
assign img[13475] = 64;
assign img[13476] = 72;
assign img[13477] = 64;
assign img[13478] = 64;
assign img[13479] = 66;
assign img[13480] = 64;
assign img[13481] = 68;
assign img[13482] = 58;
assign img[13483] = 68;
assign img[13484] = 64;
assign img[13485] = 66;
assign img[13486] = 68;
assign img[13487] = 65;
assign img[13488] = 64;
assign img[13489] = 68;
assign img[13490] = 64;
assign img[13491] = 64;
assign img[13492] = 66;
assign img[13493] = 66;
assign img[13494] = 64;
assign img[13495] = 66;
assign img[13496] = 64;
assign img[13497] = 64;
assign img[13498] = 64;
assign img[13499] = 64;
assign img[13500] = 64;
assign img[13501] = 64;
assign img[13502] = 64;
assign img[13503] = 70;
assign img[13504] = 64;
assign img[13505] = 64;
assign img[13506] = 64;
assign img[13507] = 64;
assign img[13508] = 64;
assign img[13509] = 64;
assign img[13510] = 68;
assign img[13511] = 64;
assign img[13512] = 68;
assign img[13513] = 64;
assign img[13514] = 64;
assign img[13515] = 64;
assign img[13516] = 69;
assign img[13517] = 65;
assign img[13518] = 64;
assign img[13519] = 64;
assign img[13520] = 64;
assign img[13521] = 64;
assign img[13522] = 65;
assign img[13523] = 64;
assign img[13524] = 64;
assign img[13525] = 65;
assign img[13526] = 64;
assign img[13527] = 64;
assign img[13528] = 56;
assign img[13529] = 52;
assign img[13530] = 52;
assign img[13531] = 51;
assign img[13532] = 52;
assign img[13533] = 48;
assign img[13534] = 52;
assign img[13535] = 50;
assign img[13536] = 48;
assign img[13537] = 51;
assign img[13538] = 48;
assign img[13539] = 50;
assign img[13540] = 48;
assign img[13541] = 52;
assign img[13542] = 53;
assign img[13543] = 43;
assign img[13544] = 44;
assign img[13545] = 48;
assign img[13546] = 47;
assign img[13547] = 46;
assign img[13548] = 44;
assign img[13549] = 42;
assign img[13550] = 38;
assign img[13551] = 48;
assign img[13552] = 45;
assign img[13553] = 46;
assign img[13554] = 46;
assign img[13555] = 48;
assign img[13556] = 45;
assign img[13557] = 42;
assign img[13558] = 38;
assign img[13559] = 45;
assign img[13560] = 40;
assign img[13561] = 42;
assign img[13562] = 46;
assign img[13563] = 42;
assign img[13564] = 47;
assign img[13565] = 38;
assign img[13566] = 46;
assign img[13567] = 43;
assign img[13568] = 41;
assign img[13569] = 54;
assign img[13570] = 50;
assign img[13571] = 52;
assign img[13572] = 57;
assign img[13573] = 54;
assign img[13574] = 56;
assign img[13575] = 52;
assign img[13576] = 54;
assign img[13577] = 64;
assign img[13578] = 65;
assign img[13579] = 69;
assign img[13580] = 64;
assign img[13581] = 64;
assign img[13582] = 51;
assign img[13583] = 64;
assign img[13584] = 68;
assign img[13585] = 64;
assign img[13586] = 64;
assign img[13587] = 64;
assign img[13588] = 65;
assign img[13589] = 64;
assign img[13590] = 64;
assign img[13591] = 64;
assign img[13592] = 64;
assign img[13593] = 67;
assign img[13594] = 64;
assign img[13595] = 68;
assign img[13596] = 56;
assign img[13597] = 64;
assign img[13598] = 64;
assign img[13599] = 65;
assign img[13600] = 68;
assign img[13601] = 65;
assign img[13602] = 64;
assign img[13603] = 64;
assign img[13604] = 65;
assign img[13605] = 65;
assign img[13606] = 64;
assign img[13607] = 64;
assign img[13608] = 64;
assign img[13609] = 65;
assign img[13610] = 64;
assign img[13611] = 68;
assign img[13612] = 64;
assign img[13613] = 55;
assign img[13614] = 66;
assign img[13615] = 67;
assign img[13616] = 69;
assign img[13617] = 68;
assign img[13618] = 64;
assign img[13619] = 64;
assign img[13620] = 57;
assign img[13621] = 64;
assign img[13622] = 65;
assign img[13623] = 64;
assign img[13624] = 65;
assign img[13625] = 65;
assign img[13626] = 64;
assign img[13627] = 64;
assign img[13628] = 65;
assign img[13629] = 64;
assign img[13630] = 66;
assign img[13631] = 68;
assign img[13632] = 65;
assign img[13633] = 65;
assign img[13634] = 64;
assign img[13635] = 65;
assign img[13636] = 57;
assign img[13637] = 64;
assign img[13638] = 66;
assign img[13639] = 64;
assign img[13640] = 54;
assign img[13641] = 65;
assign img[13642] = 65;
assign img[13643] = 57;
assign img[13644] = 66;
assign img[13645] = 64;
assign img[13646] = 64;
assign img[13647] = 64;
assign img[13648] = 59;
assign img[13649] = 58;
assign img[13650] = 61;
assign img[13651] = 64;
assign img[13652] = 66;
assign img[13653] = 57;
assign img[13654] = 64;
assign img[13655] = 64;
assign img[13656] = 57;
assign img[13657] = 48;
assign img[13658] = 46;
assign img[13659] = 44;
assign img[13660] = 42;
assign img[13661] = 50;
assign img[13662] = 44;
assign img[13663] = 41;
assign img[13664] = 41;
assign img[13665] = 46;
assign img[13666] = 40;
assign img[13667] = 43;
assign img[13668] = 45;
assign img[13669] = 44;
assign img[13670] = 39;
assign img[13671] = 48;
assign img[13672] = 43;
assign img[13673] = 43;
assign img[13674] = 44;
assign img[13675] = 41;
assign img[13676] = 39;
assign img[13677] = 47;
assign img[13678] = 40;
assign img[13679] = 38;
assign img[13680] = 45;
assign img[13681] = 42;
assign img[13682] = 41;
assign img[13683] = 41;
assign img[13684] = 46;
assign img[13685] = 38;
assign img[13686] = 40;
assign img[13687] = 36;
assign img[13688] = 36;
assign img[13689] = 37;
assign img[13690] = 40;
assign img[13691] = 37;
assign img[13692] = 34;
assign img[13693] = 41;
assign img[13694] = 37;
assign img[13695] = 37;
assign img[13696] = 32;
assign img[13697] = 65;
assign img[13698] = 66;
assign img[13699] = 70;
assign img[13700] = 68;
assign img[13701] = 64;
assign img[13702] = 67;
assign img[13703] = 67;
assign img[13704] = 68;
assign img[13705] = 72;
assign img[13706] = 72;
assign img[13707] = 73;
assign img[13708] = 81;
assign img[13709] = 76;
assign img[13710] = 73;
assign img[13711] = 75;
assign img[13712] = 69;
assign img[13713] = 77;
assign img[13714] = 75;
assign img[13715] = 80;
assign img[13716] = 73;
assign img[13717] = 73;
assign img[13718] = 73;
assign img[13719] = 82;
assign img[13720] = 79;
assign img[13721] = 80;
assign img[13722] = 82;
assign img[13723] = 80;
assign img[13724] = 77;
assign img[13725] = 69;
assign img[13726] = 77;
assign img[13727] = 81;
assign img[13728] = 76;
assign img[13729] = 81;
assign img[13730] = 73;
assign img[13731] = 81;
assign img[13732] = 75;
assign img[13733] = 76;
assign img[13734] = 81;
assign img[13735] = 77;
assign img[13736] = 75;
assign img[13737] = 81;
assign img[13738] = 73;
assign img[13739] = 78;
assign img[13740] = 75;
assign img[13741] = 72;
assign img[13742] = 85;
assign img[13743] = 78;
assign img[13744] = 77;
assign img[13745] = 77;
assign img[13746] = 72;
assign img[13747] = 80;
assign img[13748] = 73;
assign img[13749] = 77;
assign img[13750] = 70;
assign img[13751] = 74;
assign img[13752] = 77;
assign img[13753] = 78;
assign img[13754] = 80;
assign img[13755] = 81;
assign img[13756] = 73;
assign img[13757] = 81;
assign img[13758] = 84;
assign img[13759] = 77;
assign img[13760] = 77;
assign img[13761] = 77;
assign img[13762] = 76;
assign img[13763] = 74;
assign img[13764] = 79;
assign img[13765] = 77;
assign img[13766] = 79;
assign img[13767] = 77;
assign img[13768] = 76;
assign img[13769] = 70;
assign img[13770] = 76;
assign img[13771] = 76;
assign img[13772] = 76;
assign img[13773] = 76;
assign img[13774] = 72;
assign img[13775] = 78;
assign img[13776] = 75;
assign img[13777] = 78;
assign img[13778] = 76;
assign img[13779] = 82;
assign img[13780] = 78;
assign img[13781] = 76;
assign img[13782] = 76;
assign img[13783] = 65;
assign img[13784] = 66;
assign img[13785] = 64;
assign img[13786] = 64;
assign img[13787] = 64;
assign img[13788] = 64;
assign img[13789] = 64;
assign img[13790] = 64;
assign img[13791] = 64;
assign img[13792] = 64;
assign img[13793] = 64;
assign img[13794] = 64;
assign img[13795] = 64;
assign img[13796] = 54;
assign img[13797] = 64;
assign img[13798] = 64;
assign img[13799] = 64;
assign img[13800] = 64;
assign img[13801] = 64;
assign img[13802] = 54;
assign img[13803] = 64;
assign img[13804] = 65;
assign img[13805] = 64;
assign img[13806] = 54;
assign img[13807] = 64;
assign img[13808] = 64;
assign img[13809] = 52;
assign img[13810] = 64;
assign img[13811] = 51;
assign img[13812] = 46;
assign img[13813] = 51;
assign img[13814] = 53;
assign img[13815] = 53;
assign img[13816] = 64;
assign img[13817] = 46;
assign img[13818] = 52;
assign img[13819] = 49;
assign img[13820] = 54;
assign img[13821] = 53;
assign img[13822] = 64;
assign img[13823] = 64;
assign img[13824] = 52;
assign img[13825] = 69;
assign img[13826] = 67;
assign img[13827] = 68;
assign img[13828] = 70;
assign img[13829] = 73;
assign img[13830] = 72;
assign img[13831] = 75;
assign img[13832] = 73;
assign img[13833] = 64;
assign img[13834] = 74;
assign img[13835] = 88;
assign img[13836] = 81;
assign img[13837] = 80;
assign img[13838] = 80;
assign img[13839] = 77;
assign img[13840] = 81;
assign img[13841] = 80;
assign img[13842] = 82;
assign img[13843] = 84;
assign img[13844] = 81;
assign img[13845] = 82;
assign img[13846] = 84;
assign img[13847] = 81;
assign img[13848] = 76;
assign img[13849] = 84;
assign img[13850] = 83;
assign img[13851] = 85;
assign img[13852] = 82;
assign img[13853] = 82;
assign img[13854] = 82;
assign img[13855] = 85;
assign img[13856] = 86;
assign img[13857] = 80;
assign img[13858] = 81;
assign img[13859] = 84;
assign img[13860] = 81;
assign img[13861] = 81;
assign img[13862] = 81;
assign img[13863] = 79;
assign img[13864] = 88;
assign img[13865] = 85;
assign img[13866] = 82;
assign img[13867] = 86;
assign img[13868] = 97;
assign img[13869] = 85;
assign img[13870] = 84;
assign img[13871] = 85;
assign img[13872] = 89;
assign img[13873] = 88;
assign img[13874] = 84;
assign img[13875] = 77;
assign img[13876] = 85;
assign img[13877] = 85;
assign img[13878] = 86;
assign img[13879] = 88;
assign img[13880] = 82;
assign img[13881] = 84;
assign img[13882] = 82;
assign img[13883] = 84;
assign img[13884] = 85;
assign img[13885] = 82;
assign img[13886] = 78;
assign img[13887] = 90;
assign img[13888] = 81;
assign img[13889] = 85;
assign img[13890] = 90;
assign img[13891] = 88;
assign img[13892] = 83;
assign img[13893] = 83;
assign img[13894] = 80;
assign img[13895] = 84;
assign img[13896] = 76;
assign img[13897] = 80;
assign img[13898] = 87;
assign img[13899] = 81;
assign img[13900] = 82;
assign img[13901] = 81;
assign img[13902] = 82;
assign img[13903] = 82;
assign img[13904] = 79;
assign img[13905] = 80;
assign img[13906] = 84;
assign img[13907] = 86;
assign img[13908] = 80;
assign img[13909] = 83;
assign img[13910] = 80;
assign img[13911] = 78;
assign img[13912] = 72;
assign img[13913] = 72;
assign img[13914] = 64;
assign img[13915] = 71;
assign img[13916] = 70;
assign img[13917] = 74;
assign img[13918] = 64;
assign img[13919] = 68;
assign img[13920] = 70;
assign img[13921] = 68;
assign img[13922] = 64;
assign img[13923] = 65;
assign img[13924] = 66;
assign img[13925] = 66;
assign img[13926] = 64;
assign img[13927] = 64;
assign img[13928] = 64;
assign img[13929] = 64;
assign img[13930] = 64;
assign img[13931] = 64;
assign img[13932] = 64;
assign img[13933] = 64;
assign img[13934] = 66;
assign img[13935] = 64;
assign img[13936] = 64;
assign img[13937] = 64;
assign img[13938] = 64;
assign img[13939] = 66;
assign img[13940] = 64;
assign img[13941] = 64;
assign img[13942] = 64;
assign img[13943] = 56;
assign img[13944] = 60;
assign img[13945] = 64;
assign img[13946] = 57;
assign img[13947] = 54;
assign img[13948] = 64;
assign img[13949] = 64;
assign img[13950] = 64;
assign img[13951] = 60;
assign img[13952] = 64;
assign img[13953] = 75;
assign img[13954] = 68;
assign img[13955] = 66;
assign img[13956] = 66;
assign img[13957] = 68;
assign img[13958] = 72;
assign img[13959] = 78;
assign img[13960] = 80;
assign img[13961] = 75;
assign img[13962] = 73;
assign img[13963] = 79;
assign img[13964] = 80;
assign img[13965] = 79;
assign img[13966] = 74;
assign img[13967] = 86;
assign img[13968] = 80;
assign img[13969] = 91;
assign img[13970] = 84;
assign img[13971] = 81;
assign img[13972] = 84;
assign img[13973] = 84;
assign img[13974] = 85;
assign img[13975] = 87;
assign img[13976] = 88;
assign img[13977] = 85;
assign img[13978] = 85;
assign img[13979] = 82;
assign img[13980] = 85;
assign img[13981] = 81;
assign img[13982] = 81;
assign img[13983] = 85;
assign img[13984] = 81;
assign img[13985] = 84;
assign img[13986] = 96;
assign img[13987] = 89;
assign img[13988] = 81;
assign img[13989] = 89;
assign img[13990] = 78;
assign img[13991] = 86;
assign img[13992] = 81;
assign img[13993] = 85;
assign img[13994] = 86;
assign img[13995] = 82;
assign img[13996] = 88;
assign img[13997] = 81;
assign img[13998] = 83;
assign img[13999] = 87;
assign img[14000] = 81;
assign img[14001] = 82;
assign img[14002] = 82;
assign img[14003] = 84;
assign img[14004] = 84;
assign img[14005] = 84;
assign img[14006] = 81;
assign img[14007] = 81;
assign img[14008] = 81;
assign img[14009] = 83;
assign img[14010] = 77;
assign img[14011] = 90;
assign img[14012] = 85;
assign img[14013] = 84;
assign img[14014] = 85;
assign img[14015] = 81;
assign img[14016] = 81;
assign img[14017] = 81;
assign img[14018] = 83;
assign img[14019] = 81;
assign img[14020] = 81;
assign img[14021] = 85;
assign img[14022] = 88;
assign img[14023] = 89;
assign img[14024] = 80;
assign img[14025] = 81;
assign img[14026] = 81;
assign img[14027] = 80;
assign img[14028] = 81;
assign img[14029] = 80;
assign img[14030] = 84;
assign img[14031] = 82;
assign img[14032] = 78;
assign img[14033] = 88;
assign img[14034] = 75;
assign img[14035] = 82;
assign img[14036] = 87;
assign img[14037] = 80;
assign img[14038] = 79;
assign img[14039] = 72;
assign img[14040] = 70;
assign img[14041] = 71;
assign img[14042] = 70;
assign img[14043] = 70;
assign img[14044] = 70;
assign img[14045] = 65;
assign img[14046] = 68;
assign img[14047] = 64;
assign img[14048] = 66;
assign img[14049] = 64;
assign img[14050] = 65;
assign img[14051] = 64;
assign img[14052] = 68;
assign img[14053] = 64;
assign img[14054] = 64;
assign img[14055] = 64;
assign img[14056] = 64;
assign img[14057] = 57;
assign img[14058] = 64;
assign img[14059] = 65;
assign img[14060] = 56;
assign img[14061] = 64;
assign img[14062] = 64;
assign img[14063] = 65;
assign img[14064] = 64;
assign img[14065] = 52;
assign img[14066] = 64;
assign img[14067] = 64;
assign img[14068] = 64;
assign img[14069] = 57;
assign img[14070] = 54;
assign img[14071] = 56;
assign img[14072] = 64;
assign img[14073] = 56;
assign img[14074] = 57;
assign img[14075] = 50;
assign img[14076] = 54;
assign img[14077] = 56;
assign img[14078] = 55;
assign img[14079] = 65;
assign img[14080] = 57;
assign img[14081] = 48;
assign img[14082] = 43;
assign img[14083] = 48;
assign img[14084] = 54;
assign img[14085] = 52;
assign img[14086] = 52;
assign img[14087] = 57;
assign img[14088] = 64;
assign img[14089] = 64;
assign img[14090] = 64;
assign img[14091] = 64;
assign img[14092] = 64;
assign img[14093] = 55;
assign img[14094] = 54;
assign img[14095] = 64;
assign img[14096] = 65;
assign img[14097] = 57;
assign img[14098] = 64;
assign img[14099] = 57;
assign img[14100] = 65;
assign img[14101] = 64;
assign img[14102] = 57;
assign img[14103] = 64;
assign img[14104] = 64;
assign img[14105] = 53;
assign img[14106] = 64;
assign img[14107] = 64;
assign img[14108] = 64;
assign img[14109] = 55;
assign img[14110] = 64;
assign img[14111] = 56;
assign img[14112] = 65;
assign img[14113] = 57;
assign img[14114] = 64;
assign img[14115] = 53;
assign img[14116] = 64;
assign img[14117] = 57;
assign img[14118] = 55;
assign img[14119] = 64;
assign img[14120] = 64;
assign img[14121] = 64;
assign img[14122] = 64;
assign img[14123] = 64;
assign img[14124] = 65;
assign img[14125] = 53;
assign img[14126] = 55;
assign img[14127] = 64;
assign img[14128] = 64;
assign img[14129] = 65;
assign img[14130] = 64;
assign img[14131] = 64;
assign img[14132] = 57;
assign img[14133] = 57;
assign img[14134] = 64;
assign img[14135] = 64;
assign img[14136] = 64;
assign img[14137] = 65;
assign img[14138] = 64;
assign img[14139] = 64;
assign img[14140] = 64;
assign img[14141] = 64;
assign img[14142] = 64;
assign img[14143] = 64;
assign img[14144] = 65;
assign img[14145] = 64;
assign img[14146] = 64;
assign img[14147] = 53;
assign img[14148] = 64;
assign img[14149] = 65;
assign img[14150] = 53;
assign img[14151] = 56;
assign img[14152] = 65;
assign img[14153] = 64;
assign img[14154] = 57;
assign img[14155] = 64;
assign img[14156] = 64;
assign img[14157] = 53;
assign img[14158] = 64;
assign img[14159] = 64;
assign img[14160] = 64;
assign img[14161] = 60;
assign img[14162] = 56;
assign img[14163] = 68;
assign img[14164] = 57;
assign img[14165] = 56;
assign img[14166] = 53;
assign img[14167] = 53;
assign img[14168] = 47;
assign img[14169] = 55;
assign img[14170] = 47;
assign img[14171] = 44;
assign img[14172] = 46;
assign img[14173] = 46;
assign img[14174] = 45;
assign img[14175] = 41;
assign img[14176] = 40;
assign img[14177] = 46;
assign img[14178] = 42;
assign img[14179] = 44;
assign img[14180] = 44;
assign img[14181] = 44;
assign img[14182] = 40;
assign img[14183] = 40;
assign img[14184] = 37;
assign img[14185] = 38;
assign img[14186] = 36;
assign img[14187] = 39;
assign img[14188] = 42;
assign img[14189] = 38;
assign img[14190] = 34;
assign img[14191] = 39;
assign img[14192] = 42;
assign img[14193] = 36;
assign img[14194] = 38;
assign img[14195] = 36;
assign img[14196] = 39;
assign img[14197] = 37;
assign img[14198] = 38;
assign img[14199] = 36;
assign img[14200] = 36;
assign img[14201] = 36;
assign img[14202] = 37;
assign img[14203] = 36;
assign img[14204] = 35;
assign img[14205] = 38;
assign img[14206] = 33;
assign img[14207] = 34;
assign img[14208] = 34;
assign img[14209] = 68;
assign img[14210] = 71;
assign img[14211] = 64;
assign img[14212] = 65;
assign img[14213] = 69;
assign img[14214] = 68;
assign img[14215] = 75;
assign img[14216] = 70;
assign img[14217] = 82;
assign img[14218] = 82;
assign img[14219] = 81;
assign img[14220] = 81;
assign img[14221] = 81;
assign img[14222] = 81;
assign img[14223] = 77;
assign img[14224] = 81;
assign img[14225] = 81;
assign img[14226] = 76;
assign img[14227] = 81;
assign img[14228] = 81;
assign img[14229] = 77;
assign img[14230] = 81;
assign img[14231] = 81;
assign img[14232] = 85;
assign img[14233] = 80;
assign img[14234] = 75;
assign img[14235] = 80;
assign img[14236] = 76;
assign img[14237] = 77;
assign img[14238] = 79;
assign img[14239] = 75;
assign img[14240] = 81;
assign img[14241] = 81;
assign img[14242] = 73;
assign img[14243] = 81;
assign img[14244] = 81;
assign img[14245] = 81;
assign img[14246] = 77;
assign img[14247] = 73;
assign img[14248] = 77;
assign img[14249] = 82;
assign img[14250] = 77;
assign img[14251] = 80;
assign img[14252] = 80;
assign img[14253] = 81;
assign img[14254] = 82;
assign img[14255] = 81;
assign img[14256] = 77;
assign img[14257] = 83;
assign img[14258] = 78;
assign img[14259] = 74;
assign img[14260] = 73;
assign img[14261] = 81;
assign img[14262] = 77;
assign img[14263] = 82;
assign img[14264] = 75;
assign img[14265] = 81;
assign img[14266] = 81;
assign img[14267] = 88;
assign img[14268] = 90;
assign img[14269] = 82;
assign img[14270] = 81;
assign img[14271] = 80;
assign img[14272] = 77;
assign img[14273] = 84;
assign img[14274] = 83;
assign img[14275] = 89;
assign img[14276] = 85;
assign img[14277] = 84;
assign img[14278] = 80;
assign img[14279] = 80;
assign img[14280] = 77;
assign img[14281] = 80;
assign img[14282] = 81;
assign img[14283] = 77;
assign img[14284] = 77;
assign img[14285] = 79;
assign img[14286] = 82;
assign img[14287] = 85;
assign img[14288] = 73;
assign img[14289] = 76;
assign img[14290] = 76;
assign img[14291] = 78;
assign img[14292] = 82;
assign img[14293] = 76;
assign img[14294] = 81;
assign img[14295] = 80;
assign img[14296] = 67;
assign img[14297] = 69;
assign img[14298] = 70;
assign img[14299] = 68;
assign img[14300] = 67;
assign img[14301] = 65;
assign img[14302] = 68;
assign img[14303] = 64;
assign img[14304] = 69;
assign img[14305] = 65;
assign img[14306] = 65;
assign img[14307] = 64;
assign img[14308] = 57;
assign img[14309] = 64;
assign img[14310] = 64;
assign img[14311] = 64;
assign img[14312] = 65;
assign img[14313] = 64;
assign img[14314] = 64;
assign img[14315] = 67;
assign img[14316] = 64;
assign img[14317] = 64;
assign img[14318] = 64;
assign img[14319] = 64;
assign img[14320] = 64;
assign img[14321] = 64;
assign img[14322] = 64;
assign img[14323] = 53;
assign img[14324] = 64;
assign img[14325] = 55;
assign img[14326] = 64;
assign img[14327] = 64;
assign img[14328] = 64;
assign img[14329] = 57;
assign img[14330] = 54;
assign img[14331] = 58;
assign img[14332] = 57;
assign img[14333] = 56;
assign img[14334] = 52;
assign img[14335] = 57;
assign img[14336] = 128;
assign img[14337] = 73;
assign img[14338] = 64;
assign img[14339] = 70;
assign img[14340] = 78;
assign img[14341] = 76;
assign img[14342] = 78;
assign img[14343] = 78;
assign img[14344] = 72;
assign img[14345] = 80;
assign img[14346] = 88;
assign img[14347] = 88;
assign img[14348] = 88;
assign img[14349] = 91;
assign img[14350] = 83;
assign img[14351] = 98;
assign img[14352] = 90;
assign img[14353] = 90;
assign img[14354] = 84;
assign img[14355] = 90;
assign img[14356] = 88;
assign img[14357] = 91;
assign img[14358] = 90;
assign img[14359] = 92;
assign img[14360] = 86;
assign img[14361] = 96;
assign img[14362] = 90;
assign img[14363] = 92;
assign img[14364] = 86;
assign img[14365] = 79;
assign img[14366] = 84;
assign img[14367] = 96;
assign img[14368] = 80;
assign img[14369] = 96;
assign img[14370] = 91;
assign img[14371] = 92;
assign img[14372] = 88;
assign img[14373] = 82;
assign img[14374] = 84;
assign img[14375] = 96;
assign img[14376] = 84;
assign img[14377] = 84;
assign img[14378] = 90;
assign img[14379] = 87;
assign img[14380] = 96;
assign img[14381] = 84;
assign img[14382] = 82;
assign img[14383] = 88;
assign img[14384] = 86;
assign img[14385] = 108;
assign img[14386] = 88;
assign img[14387] = 94;
assign img[14388] = 96;
assign img[14389] = 92;
assign img[14390] = 89;
assign img[14391] = 83;
assign img[14392] = 87;
assign img[14393] = 92;
assign img[14394] = 96;
assign img[14395] = 91;
assign img[14396] = 85;
assign img[14397] = 88;
assign img[14398] = 98;
assign img[14399] = 80;
assign img[14400] = 85;
assign img[14401] = 90;
assign img[14402] = 96;
assign img[14403] = 86;
assign img[14404] = 86;
assign img[14405] = 88;
assign img[14406] = 84;
assign img[14407] = 86;
assign img[14408] = 92;
assign img[14409] = 80;
assign img[14410] = 86;
assign img[14411] = 90;
assign img[14412] = 86;
assign img[14413] = 80;
assign img[14414] = 85;
assign img[14415] = 96;
assign img[14416] = 86;
assign img[14417] = 86;
assign img[14418] = 86;
assign img[14419] = 88;
assign img[14420] = 85;
assign img[14421] = 86;
assign img[14422] = 80;
assign img[14423] = 79;
assign img[14424] = 70;
assign img[14425] = 74;
assign img[14426] = 76;
assign img[14427] = 71;
assign img[14428] = 64;
assign img[14429] = 68;
assign img[14430] = 68;
assign img[14431] = 70;
assign img[14432] = 65;
assign img[14433] = 70;
assign img[14434] = 68;
assign img[14435] = 68;
assign img[14436] = 64;
assign img[14437] = 64;
assign img[14438] = 64;
assign img[14439] = 64;
assign img[14440] = 66;
assign img[14441] = 64;
assign img[14442] = 68;
assign img[14443] = 64;
assign img[14444] = 68;
assign img[14445] = 64;
assign img[14446] = 64;
assign img[14447] = 64;
assign img[14448] = 64;
assign img[14449] = 66;
assign img[14450] = 64;
assign img[14451] = 64;
assign img[14452] = 64;
assign img[14453] = 64;
assign img[14454] = 64;
assign img[14455] = 54;
assign img[14456] = 64;
assign img[14457] = 64;
assign img[14458] = 64;
assign img[14459] = 64;
assign img[14460] = 64;
assign img[14461] = 54;
assign img[14462] = 64;
assign img[14463] = 64;
assign img[14464] = 68;
assign img[14465] = 75;
assign img[14466] = 79;
assign img[14467] = 74;
assign img[14468] = 74;
assign img[14469] = 82;
assign img[14470] = 78;
assign img[14471] = 84;
assign img[14472] = 77;
assign img[14473] = 84;
assign img[14474] = 88;
assign img[14475] = 92;
assign img[14476] = 100;
assign img[14477] = 86;
assign img[14478] = 86;
assign img[14479] = 89;
assign img[14480] = 98;
assign img[14481] = 94;
assign img[14482] = 96;
assign img[14483] = 96;
assign img[14484] = 88;
assign img[14485] = 96;
assign img[14486] = 99;
assign img[14487] = 98;
assign img[14488] = 96;
assign img[14489] = 96;
assign img[14490] = 94;
assign img[14491] = 88;
assign img[14492] = 98;
assign img[14493] = 100;
assign img[14494] = 100;
assign img[14495] = 96;
assign img[14496] = 102;
assign img[14497] = 102;
assign img[14498] = 96;
assign img[14499] = 100;
assign img[14500] = 88;
assign img[14501] = 87;
assign img[14502] = 96;
assign img[14503] = 97;
assign img[14504] = 94;
assign img[14505] = 102;
assign img[14506] = 102;
assign img[14507] = 95;
assign img[14508] = 102;
assign img[14509] = 87;
assign img[14510] = 102;
assign img[14511] = 94;
assign img[14512] = 98;
assign img[14513] = 98;
assign img[14514] = 96;
assign img[14515] = 98;
assign img[14516] = 98;
assign img[14517] = 94;
assign img[14518] = 102;
assign img[14519] = 94;
assign img[14520] = 92;
assign img[14521] = 95;
assign img[14522] = 92;
assign img[14523] = 90;
assign img[14524] = 92;
assign img[14525] = 88;
assign img[14526] = 89;
assign img[14527] = 89;
assign img[14528] = 96;
assign img[14529] = 96;
assign img[14530] = 84;
assign img[14531] = 86;
assign img[14532] = 87;
assign img[14533] = 96;
assign img[14534] = 96;
assign img[14535] = 88;
assign img[14536] = 88;
assign img[14537] = 92;
assign img[14538] = 88;
assign img[14539] = 92;
assign img[14540] = 80;
assign img[14541] = 92;
assign img[14542] = 96;
assign img[14543] = 86;
assign img[14544] = 96;
assign img[14545] = 99;
assign img[14546] = 92;
assign img[14547] = 92;
assign img[14548] = 80;
assign img[14549] = 86;
assign img[14550] = 84;
assign img[14551] = 80;
assign img[14552] = 80;
assign img[14553] = 87;
assign img[14554] = 79;
assign img[14555] = 72;
assign img[14556] = 78;
assign img[14557] = 76;
assign img[14558] = 72;
assign img[14559] = 73;
assign img[14560] = 72;
assign img[14561] = 76;
assign img[14562] = 71;
assign img[14563] = 72;
assign img[14564] = 71;
assign img[14565] = 76;
assign img[14566] = 69;
assign img[14567] = 68;
assign img[14568] = 68;
assign img[14569] = 68;
assign img[14570] = 72;
assign img[14571] = 68;
assign img[14572] = 68;
assign img[14573] = 77;
assign img[14574] = 72;
assign img[14575] = 68;
assign img[14576] = 68;
assign img[14577] = 72;
assign img[14578] = 64;
assign img[14579] = 64;
assign img[14580] = 64;
assign img[14581] = 64;
assign img[14582] = 65;
assign img[14583] = 64;
assign img[14584] = 64;
assign img[14585] = 76;
assign img[14586] = 65;
assign img[14587] = 68;
assign img[14588] = 68;
assign img[14589] = 60;
assign img[14590] = 68;
assign img[14591] = 65;
assign img[14592] = 68;
assign img[14593] = 96;
assign img[14594] = 95;
assign img[14595] = 96;
assign img[14596] = 108;
assign img[14597] = 100;
assign img[14598] = 111;
assign img[14599] = 128;
assign img[14600] = 104;
assign img[14601] = 128;
assign img[14602] = 128;
assign img[14603] = 128;
assign img[14604] = 128;
assign img[14605] = 128;
assign img[14606] = 111;
assign img[14607] = 128;
assign img[14608] = 128;
assign img[14609] = 128;
assign img[14610] = 112;
assign img[14611] = 128;
assign img[14612] = 128;
assign img[14613] = 128;
assign img[14614] = 128;
assign img[14615] = 128;
assign img[14616] = 112;
assign img[14617] = 128;
assign img[14618] = 128;
assign img[14619] = 128;
assign img[14620] = 128;
assign img[14621] = 128;
assign img[14622] = 128;
assign img[14623] = 128;
assign img[14624] = 128;
assign img[14625] = 128;
assign img[14626] = 128;
assign img[14627] = 128;
assign img[14628] = 110;
assign img[14629] = 128;
assign img[14630] = 128;
assign img[14631] = 128;
assign img[14632] = 128;
assign img[14633] = 128;
assign img[14634] = 112;
assign img[14635] = 128;
assign img[14636] = 128;
assign img[14637] = 128;
assign img[14638] = 128;
assign img[14639] = 128;
assign img[14640] = 128;
assign img[14641] = 128;
assign img[14642] = 114;
assign img[14643] = 118;
assign img[14644] = 128;
assign img[14645] = 129;
assign img[14646] = 128;
assign img[14647] = 128;
assign img[14648] = 128;
assign img[14649] = 128;
assign img[14650] = 128;
assign img[14651] = 128;
assign img[14652] = 128;
assign img[14653] = 128;
assign img[14654] = 128;
assign img[14655] = 128;
assign img[14656] = 128;
assign img[14657] = 128;
assign img[14658] = 128;
assign img[14659] = 128;
assign img[14660] = 112;
assign img[14661] = 128;
assign img[14662] = 128;
assign img[14663] = 109;
assign img[14664] = 128;
assign img[14665] = 128;
assign img[14666] = 128;
assign img[14667] = 128;
assign img[14668] = 128;
assign img[14669] = 128;
assign img[14670] = 128;
assign img[14671] = 128;
assign img[14672] = 111;
assign img[14673] = 128;
assign img[14674] = 128;
assign img[14675] = 128;
assign img[14676] = 116;
assign img[14677] = 128;
assign img[14678] = 128;
assign img[14679] = 111;
assign img[14680] = 104;
assign img[14681] = 105;
assign img[14682] = 128;
assign img[14683] = 108;
assign img[14684] = 100;
assign img[14685] = 92;
assign img[14686] = 95;
assign img[14687] = 94;
assign img[14688] = 93;
assign img[14689] = 100;
assign img[14690] = 99;
assign img[14691] = 92;
assign img[14692] = 92;
assign img[14693] = 96;
assign img[14694] = 86;
assign img[14695] = 102;
assign img[14696] = 92;
assign img[14697] = 89;
assign img[14698] = 95;
assign img[14699] = 96;
assign img[14700] = 89;
assign img[14701] = 92;
assign img[14702] = 96;
assign img[14703] = 95;
assign img[14704] = 92;
assign img[14705] = 96;
assign img[14706] = 89;
assign img[14707] = 92;
assign img[14708] = 92;
assign img[14709] = 94;
assign img[14710] = 80;
assign img[14711] = 88;
assign img[14712] = 92;
assign img[14713] = 81;
assign img[14714] = 84;
assign img[14715] = 85;
assign img[14716] = 96;
assign img[14717] = 93;
assign img[14718] = 96;
assign img[14719] = 84;
assign img[14720] = 80;
assign img[14721] = 88;
assign img[14722] = 92;
assign img[14723] = 90;
assign img[14724] = 94;
assign img[14725] = 97;
assign img[14726] = 98;
assign img[14727] = 102;
assign img[14728] = 102;
assign img[14729] = 112;
assign img[14730] = 114;
assign img[14731] = 112;
assign img[14732] = 111;
assign img[14733] = 110;
assign img[14734] = 128;
assign img[14735] = 112;
assign img[14736] = 110;
assign img[14737] = 128;
assign img[14738] = 128;
assign img[14739] = 111;
assign img[14740] = 111;
assign img[14741] = 111;
assign img[14742] = 128;
assign img[14743] = 128;
assign img[14744] = 112;
assign img[14745] = 110;
assign img[14746] = 111;
assign img[14747] = 110;
assign img[14748] = 111;
assign img[14749] = 111;
assign img[14750] = 110;
assign img[14751] = 128;
assign img[14752] = 128;
assign img[14753] = 112;
assign img[14754] = 111;
assign img[14755] = 111;
assign img[14756] = 128;
assign img[14757] = 104;
assign img[14758] = 111;
assign img[14759] = 111;
assign img[14760] = 111;
assign img[14761] = 108;
assign img[14762] = 112;
assign img[14763] = 111;
assign img[14764] = 112;
assign img[14765] = 111;
assign img[14766] = 111;
assign img[14767] = 128;
assign img[14768] = 110;
assign img[14769] = 104;
assign img[14770] = 110;
assign img[14771] = 108;
assign img[14772] = 110;
assign img[14773] = 106;
assign img[14774] = 102;
assign img[14775] = 114;
assign img[14776] = 112;
assign img[14777] = 112;
assign img[14778] = 111;
assign img[14779] = 111;
assign img[14780] = 110;
assign img[14781] = 108;
assign img[14782] = 105;
assign img[14783] = 128;
assign img[14784] = 105;
assign img[14785] = 104;
assign img[14786] = 101;
assign img[14787] = 104;
assign img[14788] = 111;
assign img[14789] = 105;
assign img[14790] = 128;
assign img[14791] = 100;
assign img[14792] = 108;
assign img[14793] = 110;
assign img[14794] = 128;
assign img[14795] = 107;
assign img[14796] = 128;
assign img[14797] = 128;
assign img[14798] = 105;
assign img[14799] = 104;
assign img[14800] = 110;
assign img[14801] = 113;
assign img[14802] = 107;
assign img[14803] = 105;
assign img[14804] = 108;
assign img[14805] = 104;
assign img[14806] = 98;
assign img[14807] = 108;
assign img[14808] = 98;
assign img[14809] = 90;
assign img[14810] = 90;
assign img[14811] = 94;
assign img[14812] = 91;
assign img[14813] = 93;
assign img[14814] = 94;
assign img[14815] = 95;
assign img[14816] = 88;
assign img[14817] = 92;
assign img[14818] = 86;
assign img[14819] = 90;
assign img[14820] = 92;
assign img[14821] = 89;
assign img[14822] = 96;
assign img[14823] = 89;
assign img[14824] = 96;
assign img[14825] = 84;
assign img[14826] = 94;
assign img[14827] = 80;
assign img[14828] = 80;
assign img[14829] = 82;
assign img[14830] = 81;
assign img[14831] = 80;
assign img[14832] = 84;
assign img[14833] = 82;
assign img[14834] = 78;
assign img[14835] = 84;
assign img[14836] = 84;
assign img[14837] = 84;
assign img[14838] = 79;
assign img[14839] = 85;
assign img[14840] = 80;
assign img[14841] = 80;
assign img[14842] = 84;
assign img[14843] = 88;
assign img[14844] = 80;
assign img[14845] = 76;
assign img[14846] = 76;
assign img[14847] = 82;
assign img[14848] = 80;
assign img[14849] = 73;
assign img[14850] = 68;
assign img[14851] = 74;
assign img[14852] = 75;
assign img[14853] = 81;
assign img[14854] = 76;
assign img[14855] = 81;
assign img[14856] = 77;
assign img[14857] = 80;
assign img[14858] = 88;
assign img[14859] = 96;
assign img[14860] = 86;
assign img[14861] = 84;
assign img[14862] = 90;
assign img[14863] = 86;
assign img[14864] = 92;
assign img[14865] = 86;
assign img[14866] = 86;
assign img[14867] = 96;
assign img[14868] = 86;
assign img[14869] = 86;
assign img[14870] = 96;
assign img[14871] = 88;
assign img[14872] = 86;
assign img[14873] = 96;
assign img[14874] = 88;
assign img[14875] = 89;
assign img[14876] = 96;
assign img[14877] = 86;
assign img[14878] = 86;
assign img[14879] = 88;
assign img[14880] = 90;
assign img[14881] = 95;
assign img[14882] = 92;
assign img[14883] = 92;
assign img[14884] = 98;
assign img[14885] = 88;
assign img[14886] = 92;
assign img[14887] = 86;
assign img[14888] = 96;
assign img[14889] = 88;
assign img[14890] = 87;
assign img[14891] = 98;
assign img[14892] = 87;
assign img[14893] = 84;
assign img[14894] = 92;
assign img[14895] = 96;
assign img[14896] = 88;
assign img[14897] = 98;
assign img[14898] = 98;
assign img[14899] = 98;
assign img[14900] = 92;
assign img[14901] = 90;
assign img[14902] = 90;
assign img[14903] = 96;
assign img[14904] = 92;
assign img[14905] = 102;
assign img[14906] = 92;
assign img[14907] = 86;
assign img[14908] = 92;
assign img[14909] = 89;
assign img[14910] = 84;
assign img[14911] = 88;
assign img[14912] = 85;
assign img[14913] = 89;
assign img[14914] = 85;
assign img[14915] = 93;
assign img[14916] = 88;
assign img[14917] = 92;
assign img[14918] = 88;
assign img[14919] = 88;
assign img[14920] = 86;
assign img[14921] = 88;
assign img[14922] = 90;
assign img[14923] = 89;
assign img[14924] = 80;
assign img[14925] = 80;
assign img[14926] = 88;
assign img[14927] = 89;
assign img[14928] = 88;
assign img[14929] = 85;
assign img[14930] = 88;
assign img[14931] = 86;
assign img[14932] = 90;
assign img[14933] = 81;
assign img[14934] = 79;
assign img[14935] = 73;
assign img[14936] = 74;
assign img[14937] = 76;
assign img[14938] = 73;
assign img[14939] = 76;
assign img[14940] = 68;
assign img[14941] = 74;
assign img[14942] = 72;
assign img[14943] = 73;
assign img[14944] = 65;
assign img[14945] = 65;
assign img[14946] = 72;
assign img[14947] = 65;
assign img[14948] = 73;
assign img[14949] = 64;
assign img[14950] = 72;
assign img[14951] = 64;
assign img[14952] = 66;
assign img[14953] = 68;
assign img[14954] = 72;
assign img[14955] = 68;
assign img[14956] = 68;
assign img[14957] = 68;
assign img[14958] = 72;
assign img[14959] = 64;
assign img[14960] = 64;
assign img[14961] = 67;
assign img[14962] = 72;
assign img[14963] = 60;
assign img[14964] = 64;
assign img[14965] = 64;
assign img[14966] = 71;
assign img[14967] = 66;
assign img[14968] = 68;
assign img[14969] = 65;
assign img[14970] = 68;
assign img[14971] = 58;
assign img[14972] = 64;
assign img[14973] = 57;
assign img[14974] = 64;
assign img[14975] = 68;
assign img[14976] = 54;
assign img[14977] = 96;
assign img[14978] = 89;
assign img[14979] = 88;
assign img[14980] = 89;
assign img[14981] = 96;
assign img[14982] = 96;
assign img[14983] = 92;
assign img[14984] = 88;
assign img[14985] = 102;
assign img[14986] = 109;
assign img[14987] = 102;
assign img[14988] = 110;
assign img[14989] = 104;
assign img[14990] = 102;
assign img[14991] = 104;
assign img[14992] = 102;
assign img[14993] = 110;
assign img[14994] = 110;
assign img[14995] = 103;
assign img[14996] = 103;
assign img[14997] = 104;
assign img[14998] = 111;
assign img[14999] = 102;
assign img[15000] = 100;
assign img[15001] = 104;
assign img[15002] = 110;
assign img[15003] = 111;
assign img[15004] = 100;
assign img[15005] = 110;
assign img[15006] = 111;
assign img[15007] = 103;
assign img[15008] = 110;
assign img[15009] = 110;
assign img[15010] = 103;
assign img[15011] = 102;
assign img[15012] = 98;
assign img[15013] = 104;
assign img[15014] = 103;
assign img[15015] = 102;
assign img[15016] = 103;
assign img[15017] = 103;
assign img[15018] = 99;
assign img[15019] = 104;
assign img[15020] = 99;
assign img[15021] = 104;
assign img[15022] = 111;
assign img[15023] = 104;
assign img[15024] = 101;
assign img[15025] = 106;
assign img[15026] = 104;
assign img[15027] = 110;
assign img[15028] = 103;
assign img[15029] = 104;
assign img[15030] = 111;
assign img[15031] = 104;
assign img[15032] = 107;
assign img[15033] = 104;
assign img[15034] = 103;
assign img[15035] = 104;
assign img[15036] = 104;
assign img[15037] = 104;
assign img[15038] = 104;
assign img[15039] = 100;
assign img[15040] = 98;
assign img[15041] = 105;
assign img[15042] = 98;
assign img[15043] = 96;
assign img[15044] = 105;
assign img[15045] = 105;
assign img[15046] = 100;
assign img[15047] = 98;
assign img[15048] = 104;
assign img[15049] = 100;
assign img[15050] = 104;
assign img[15051] = 112;
assign img[15052] = 96;
assign img[15053] = 97;
assign img[15054] = 104;
assign img[15055] = 100;
assign img[15056] = 102;
assign img[15057] = 106;
assign img[15058] = 100;
assign img[15059] = 98;
assign img[15060] = 96;
assign img[15061] = 93;
assign img[15062] = 88;
assign img[15063] = 87;
assign img[15064] = 92;
assign img[15065] = 84;
assign img[15066] = 88;
assign img[15067] = 87;
assign img[15068] = 88;
assign img[15069] = 85;
assign img[15070] = 88;
assign img[15071] = 81;
assign img[15072] = 82;
assign img[15073] = 80;
assign img[15074] = 85;
assign img[15075] = 79;
assign img[15076] = 80;
assign img[15077] = 80;
assign img[15078] = 82;
assign img[15079] = 82;
assign img[15080] = 77;
assign img[15081] = 80;
assign img[15082] = 89;
assign img[15083] = 81;
assign img[15084] = 78;
assign img[15085] = 78;
assign img[15086] = 77;
assign img[15087] = 80;
assign img[15088] = 80;
assign img[15089] = 73;
assign img[15090] = 70;
assign img[15091] = 80;
assign img[15092] = 80;
assign img[15093] = 73;
assign img[15094] = 71;
assign img[15095] = 75;
assign img[15096] = 77;
assign img[15097] = 79;
assign img[15098] = 82;
assign img[15099] = 79;
assign img[15100] = 73;
assign img[15101] = 76;
assign img[15102] = 73;
assign img[15103] = 78;
assign img[15104] = 74;
assign img[15105] = 82;
assign img[15106] = 88;
assign img[15107] = 88;
assign img[15108] = 78;
assign img[15109] = 96;
assign img[15110] = 89;
assign img[15111] = 85;
assign img[15112] = 90;
assign img[15113] = 96;
assign img[15114] = 100;
assign img[15115] = 106;
assign img[15116] = 108;
assign img[15117] = 100;
assign img[15118] = 104;
assign img[15119] = 96;
assign img[15120] = 98;
assign img[15121] = 106;
assign img[15122] = 98;
assign img[15123] = 100;
assign img[15124] = 99;
assign img[15125] = 104;
assign img[15126] = 110;
assign img[15127] = 99;
assign img[15128] = 110;
assign img[15129] = 108;
assign img[15130] = 104;
assign img[15131] = 101;
assign img[15132] = 108;
assign img[15133] = 105;
assign img[15134] = 101;
assign img[15135] = 102;
assign img[15136] = 96;
assign img[15137] = 103;
assign img[15138] = 108;
assign img[15139] = 106;
assign img[15140] = 105;
assign img[15141] = 110;
assign img[15142] = 105;
assign img[15143] = 101;
assign img[15144] = 101;
assign img[15145] = 105;
assign img[15146] = 102;
assign img[15147] = 102;
assign img[15148] = 112;
assign img[15149] = 96;
assign img[15150] = 97;
assign img[15151] = 97;
assign img[15152] = 105;
assign img[15153] = 104;
assign img[15154] = 104;
assign img[15155] = 105;
assign img[15156] = 100;
assign img[15157] = 97;
assign img[15158] = 97;
assign img[15159] = 105;
assign img[15160] = 101;
assign img[15161] = 108;
assign img[15162] = 103;
assign img[15163] = 102;
assign img[15164] = 100;
assign img[15165] = 105;
assign img[15166] = 106;
assign img[15167] = 97;
assign img[15168] = 105;
assign img[15169] = 98;
assign img[15170] = 98;
assign img[15171] = 108;
assign img[15172] = 97;
assign img[15173] = 96;
assign img[15174] = 93;
assign img[15175] = 96;
assign img[15176] = 104;
assign img[15177] = 100;
assign img[15178] = 100;
assign img[15179] = 100;
assign img[15180] = 100;
assign img[15181] = 97;
assign img[15182] = 100;
assign img[15183] = 104;
assign img[15184] = 104;
assign img[15185] = 102;
assign img[15186] = 94;
assign img[15187] = 100;
assign img[15188] = 96;
assign img[15189] = 88;
assign img[15190] = 77;
assign img[15191] = 88;
assign img[15192] = 86;
assign img[15193] = 85;
assign img[15194] = 80;
assign img[15195] = 82;
assign img[15196] = 92;
assign img[15197] = 85;
assign img[15198] = 84;
assign img[15199] = 81;
assign img[15200] = 85;
assign img[15201] = 82;
assign img[15202] = 77;
assign img[15203] = 79;
assign img[15204] = 81;
assign img[15205] = 82;
assign img[15206] = 84;
assign img[15207] = 76;
assign img[15208] = 77;
assign img[15209] = 80;
assign img[15210] = 84;
assign img[15211] = 84;
assign img[15212] = 81;
assign img[15213] = 82;
assign img[15214] = 80;
assign img[15215] = 79;
assign img[15216] = 79;
assign img[15217] = 77;
assign img[15218] = 71;
assign img[15219] = 79;
assign img[15220] = 76;
assign img[15221] = 76;
assign img[15222] = 73;
assign img[15223] = 78;
assign img[15224] = 73;
assign img[15225] = 71;
assign img[15226] = 76;
assign img[15227] = 76;
assign img[15228] = 72;
assign img[15229] = 80;
assign img[15230] = 78;
assign img[15231] = 74;
assign img[15232] = 78;
assign img[15233] = 97;
assign img[15234] = 96;
assign img[15235] = 96;
assign img[15236] = 100;
assign img[15237] = 109;
assign img[15238] = 97;
assign img[15239] = 105;
assign img[15240] = 104;
assign img[15241] = 112;
assign img[15242] = 109;
assign img[15243] = 114;
assign img[15244] = 128;
assign img[15245] = 109;
assign img[15246] = 128;
assign img[15247] = 128;
assign img[15248] = 128;
assign img[15249] = 128;
assign img[15250] = 128;
assign img[15251] = 128;
assign img[15252] = 109;
assign img[15253] = 128;
assign img[15254] = 129;
assign img[15255] = 128;
assign img[15256] = 128;
assign img[15257] = 128;
assign img[15258] = 128;
assign img[15259] = 128;
assign img[15260] = 128;
assign img[15261] = 128;
assign img[15262] = 109;
assign img[15263] = 112;
assign img[15264] = 128;
assign img[15265] = 128;
assign img[15266] = 128;
assign img[15267] = 106;
assign img[15268] = 113;
assign img[15269] = 128;
assign img[15270] = 128;
assign img[15271] = 112;
assign img[15272] = 113;
assign img[15273] = 128;
assign img[15274] = 128;
assign img[15275] = 128;
assign img[15276] = 113;
assign img[15277] = 128;
assign img[15278] = 128;
assign img[15279] = 128;
assign img[15280] = 113;
assign img[15281] = 128;
assign img[15282] = 128;
assign img[15283] = 128;
assign img[15284] = 128;
assign img[15285] = 113;
assign img[15286] = 110;
assign img[15287] = 113;
assign img[15288] = 128;
assign img[15289] = 128;
assign img[15290] = 128;
assign img[15291] = 128;
assign img[15292] = 113;
assign img[15293] = 128;
assign img[15294] = 128;
assign img[15295] = 128;
assign img[15296] = 128;
assign img[15297] = 128;
assign img[15298] = 112;
assign img[15299] = 128;
assign img[15300] = 128;
assign img[15301] = 128;
assign img[15302] = 128;
assign img[15303] = 128;
assign img[15304] = 113;
assign img[15305] = 112;
assign img[15306] = 128;
assign img[15307] = 128;
assign img[15308] = 128;
assign img[15309] = 128;
assign img[15310] = 128;
assign img[15311] = 128;
assign img[15312] = 105;
assign img[15313] = 128;
assign img[15314] = 110;
assign img[15315] = 110;
assign img[15316] = 103;
assign img[15317] = 100;
assign img[15318] = 96;
assign img[15319] = 101;
assign img[15320] = 96;
assign img[15321] = 105;
assign img[15322] = 96;
assign img[15323] = 96;
assign img[15324] = 96;
assign img[15325] = 88;
assign img[15326] = 92;
assign img[15327] = 92;
assign img[15328] = 96;
assign img[15329] = 104;
assign img[15330] = 97;
assign img[15331] = 93;
assign img[15332] = 96;
assign img[15333] = 96;
assign img[15334] = 96;
assign img[15335] = 96;
assign img[15336] = 92;
assign img[15337] = 87;
assign img[15338] = 97;
assign img[15339] = 97;
assign img[15340] = 100;
assign img[15341] = 85;
assign img[15342] = 97;
assign img[15343] = 96;
assign img[15344] = 90;
assign img[15345] = 96;
assign img[15346] = 89;
assign img[15347] = 92;
assign img[15348] = 80;
assign img[15349] = 88;
assign img[15350] = 87;
assign img[15351] = 80;
assign img[15352] = 93;
assign img[15353] = 100;
assign img[15354] = 86;
assign img[15355] = 86;
assign img[15356] = 86;
assign img[15357] = 84;
assign img[15358] = 96;
assign img[15359] = 88;
assign img[15360] = 79;
assign img[15361] = 92;
assign img[15362] = 85;
assign img[15363] = 88;
assign img[15364] = 93;
assign img[15365] = 92;
assign img[15366] = 92;
assign img[15367] = 89;
assign img[15368] = 101;
assign img[15369] = 98;
assign img[15370] = 96;
assign img[15371] = 99;
assign img[15372] = 98;
assign img[15373] = 107;
assign img[15374] = 128;
assign img[15375] = 128;
assign img[15376] = 101;
assign img[15377] = 105;
assign img[15378] = 111;
assign img[15379] = 107;
assign img[15380] = 106;
assign img[15381] = 105;
assign img[15382] = 128;
assign img[15383] = 105;
assign img[15384] = 128;
assign img[15385] = 102;
assign img[15386] = 108;
assign img[15387] = 108;
assign img[15388] = 101;
assign img[15389] = 105;
assign img[15390] = 110;
assign img[15391] = 128;
assign img[15392] = 109;
assign img[15393] = 107;
assign img[15394] = 97;
assign img[15395] = 110;
assign img[15396] = 113;
assign img[15397] = 97;
assign img[15398] = 104;
assign img[15399] = 113;
assign img[15400] = 110;
assign img[15401] = 112;
assign img[15402] = 108;
assign img[15403] = 104;
assign img[15404] = 105;
assign img[15405] = 100;
assign img[15406] = 106;
assign img[15407] = 112;
assign img[15408] = 109;
assign img[15409] = 108;
assign img[15410] = 114;
assign img[15411] = 109;
assign img[15412] = 107;
assign img[15413] = 105;
assign img[15414] = 105;
assign img[15415] = 112;
assign img[15416] = 128;
assign img[15417] = 111;
assign img[15418] = 108;
assign img[15419] = 106;
assign img[15420] = 112;
assign img[15421] = 108;
assign img[15422] = 100;
assign img[15423] = 106;
assign img[15424] = 106;
assign img[15425] = 109;
assign img[15426] = 105;
assign img[15427] = 107;
assign img[15428] = 102;
assign img[15429] = 128;
assign img[15430] = 112;
assign img[15431] = 106;
assign img[15432] = 106;
assign img[15433] = 128;
assign img[15434] = 112;
assign img[15435] = 108;
assign img[15436] = 104;
assign img[15437] = 110;
assign img[15438] = 106;
assign img[15439] = 108;
assign img[15440] = 102;
assign img[15441] = 97;
assign img[15442] = 104;
assign img[15443] = 92;
assign img[15444] = 91;
assign img[15445] = 100;
assign img[15446] = 85;
assign img[15447] = 96;
assign img[15448] = 86;
assign img[15449] = 86;
assign img[15450] = 84;
assign img[15451] = 86;
assign img[15452] = 87;
assign img[15453] = 84;
assign img[15454] = 94;
assign img[15455] = 86;
assign img[15456] = 92;
assign img[15457] = 82;
assign img[15458] = 86;
assign img[15459] = 92;
assign img[15460] = 84;
assign img[15461] = 80;
assign img[15462] = 81;
assign img[15463] = 81;
assign img[15464] = 82;
assign img[15465] = 80;
assign img[15466] = 85;
assign img[15467] = 81;
assign img[15468] = 87;
assign img[15469] = 81;
assign img[15470] = 86;
assign img[15471] = 86;
assign img[15472] = 80;
assign img[15473] = 81;
assign img[15474] = 85;
assign img[15475] = 79;
assign img[15476] = 80;
assign img[15477] = 81;
assign img[15478] = 80;
assign img[15479] = 75;
assign img[15480] = 77;
assign img[15481] = 78;
assign img[15482] = 77;
assign img[15483] = 90;
assign img[15484] = 74;
assign img[15485] = 80;
assign img[15486] = 72;
assign img[15487] = 73;
assign img[15488] = 80;
assign img[15489] = 78;
assign img[15490] = 73;
assign img[15491] = 73;
assign img[15492] = 72;
assign img[15493] = 77;
assign img[15494] = 84;
assign img[15495] = 78;
assign img[15496] = 76;
assign img[15497] = 92;
assign img[15498] = 75;
assign img[15499] = 89;
assign img[15500] = 92;
assign img[15501] = 92;
assign img[15502] = 81;
assign img[15503] = 95;
assign img[15504] = 92;
assign img[15505] = 104;
assign img[15506] = 93;
assign img[15507] = 89;
assign img[15508] = 93;
assign img[15509] = 96;
assign img[15510] = 92;
assign img[15511] = 88;
assign img[15512] = 92;
assign img[15513] = 96;
assign img[15514] = 92;
assign img[15515] = 87;
assign img[15516] = 88;
assign img[15517] = 95;
assign img[15518] = 100;
assign img[15519] = 96;
assign img[15520] = 97;
assign img[15521] = 91;
assign img[15522] = 96;
assign img[15523] = 88;
assign img[15524] = 96;
assign img[15525] = 92;
assign img[15526] = 92;
assign img[15527] = 92;
assign img[15528] = 88;
assign img[15529] = 93;
assign img[15530] = 96;
assign img[15531] = 92;
assign img[15532] = 95;
assign img[15533] = 88;
assign img[15534] = 94;
assign img[15535] = 88;
assign img[15536] = 96;
assign img[15537] = 96;
assign img[15538] = 96;
assign img[15539] = 92;
assign img[15540] = 90;
assign img[15541] = 88;
assign img[15542] = 100;
assign img[15543] = 99;
assign img[15544] = 96;
assign img[15545] = 88;
assign img[15546] = 88;
assign img[15547] = 104;
assign img[15548] = 96;
assign img[15549] = 98;
assign img[15550] = 96;
assign img[15551] = 92;
assign img[15552] = 92;
assign img[15553] = 96;
assign img[15554] = 88;
assign img[15555] = 96;
assign img[15556] = 96;
assign img[15557] = 96;
assign img[15558] = 96;
assign img[15559] = 96;
assign img[15560] = 86;
assign img[15561] = 96;
assign img[15562] = 96;
assign img[15563] = 100;
assign img[15564] = 96;
assign img[15565] = 88;
assign img[15566] = 83;
assign img[15567] = 81;
assign img[15568] = 80;
assign img[15569] = 82;
assign img[15570] = 81;
assign img[15571] = 80;
assign img[15572] = 83;
assign img[15573] = 75;
assign img[15574] = 76;
assign img[15575] = 76;
assign img[15576] = 70;
assign img[15577] = 80;
assign img[15578] = 70;
assign img[15579] = 76;
assign img[15580] = 76;
assign img[15581] = 76;
assign img[15582] = 74;
assign img[15583] = 78;
assign img[15584] = 72;
assign img[15585] = 67;
assign img[15586] = 70;
assign img[15587] = 76;
assign img[15588] = 70;
assign img[15589] = 64;
assign img[15590] = 72;
assign img[15591] = 76;
assign img[15592] = 72;
assign img[15593] = 68;
assign img[15594] = 64;
assign img[15595] = 69;
assign img[15596] = 68;
assign img[15597] = 78;
assign img[15598] = 64;
assign img[15599] = 70;
assign img[15600] = 72;
assign img[15601] = 70;
assign img[15602] = 72;
assign img[15603] = 72;
assign img[15604] = 69;
assign img[15605] = 66;
assign img[15606] = 66;
assign img[15607] = 69;
assign img[15608] = 68;
assign img[15609] = 70;
assign img[15610] = 66;
assign img[15611] = 64;
assign img[15612] = 71;
assign img[15613] = 68;
assign img[15614] = 70;
assign img[15615] = 70;
assign img[15616] = 69;
assign img[15617] = 102;
assign img[15618] = 94;
assign img[15619] = 88;
assign img[15620] = 87;
assign img[15621] = 92;
assign img[15622] = 97;
assign img[15623] = 102;
assign img[15624] = 96;
assign img[15625] = 98;
assign img[15626] = 101;
assign img[15627] = 98;
assign img[15628] = 96;
assign img[15629] = 105;
assign img[15630] = 102;
assign img[15631] = 110;
assign img[15632] = 111;
assign img[15633] = 109;
assign img[15634] = 113;
assign img[15635] = 108;
assign img[15636] = 128;
assign img[15637] = 108;
assign img[15638] = 105;
assign img[15639] = 108;
assign img[15640] = 110;
assign img[15641] = 112;
assign img[15642] = 112;
assign img[15643] = 109;
assign img[15644] = 106;
assign img[15645] = 108;
assign img[15646] = 110;
assign img[15647] = 112;
assign img[15648] = 128;
assign img[15649] = 113;
assign img[15650] = 112;
assign img[15651] = 108;
assign img[15652] = 101;
assign img[15653] = 105;
assign img[15654] = 110;
assign img[15655] = 112;
assign img[15656] = 109;
assign img[15657] = 106;
assign img[15658] = 113;
assign img[15659] = 108;
assign img[15660] = 104;
assign img[15661] = 109;
assign img[15662] = 110;
assign img[15663] = 108;
assign img[15664] = 108;
assign img[15665] = 108;
assign img[15666] = 108;
assign img[15667] = 108;
assign img[15668] = 101;
assign img[15669] = 108;
assign img[15670] = 106;
assign img[15671] = 105;
assign img[15672] = 107;
assign img[15673] = 128;
assign img[15674] = 113;
assign img[15675] = 112;
assign img[15676] = 112;
assign img[15677] = 107;
assign img[15678] = 102;
assign img[15679] = 113;
assign img[15680] = 100;
assign img[15681] = 104;
assign img[15682] = 105;
assign img[15683] = 106;
assign img[15684] = 109;
assign img[15685] = 105;
assign img[15686] = 113;
assign img[15687] = 111;
assign img[15688] = 106;
assign img[15689] = 105;
assign img[15690] = 112;
assign img[15691] = 101;
assign img[15692] = 112;
assign img[15693] = 108;
assign img[15694] = 97;
assign img[15695] = 101;
assign img[15696] = 97;
assign img[15697] = 100;
assign img[15698] = 96;
assign img[15699] = 96;
assign img[15700] = 96;
assign img[15701] = 82;
assign img[15702] = 85;
assign img[15703] = 86;
assign img[15704] = 85;
assign img[15705] = 86;
assign img[15706] = 90;
assign img[15707] = 84;
assign img[15708] = 86;
assign img[15709] = 84;
assign img[15710] = 96;
assign img[15711] = 85;
assign img[15712] = 85;
assign img[15713] = 86;
assign img[15714] = 87;
assign img[15715] = 84;
assign img[15716] = 89;
assign img[15717] = 85;
assign img[15718] = 91;
assign img[15719] = 88;
assign img[15720] = 88;
assign img[15721] = 88;
assign img[15722] = 90;
assign img[15723] = 82;
assign img[15724] = 87;
assign img[15725] = 80;
assign img[15726] = 84;
assign img[15727] = 73;
assign img[15728] = 85;
assign img[15729] = 89;
assign img[15730] = 86;
assign img[15731] = 87;
assign img[15732] = 84;
assign img[15733] = 74;
assign img[15734] = 88;
assign img[15735] = 80;
assign img[15736] = 77;
assign img[15737] = 80;
assign img[15738] = 80;
assign img[15739] = 73;
assign img[15740] = 73;
assign img[15741] = 81;
assign img[15742] = 85;
assign img[15743] = 77;
assign img[15744] = 82;
assign img[15745] = 86;
assign img[15746] = 96;
assign img[15747] = 87;
assign img[15748] = 87;
assign img[15749] = 86;
assign img[15750] = 90;
assign img[15751] = 104;
assign img[15752] = 84;
assign img[15753] = 96;
assign img[15754] = 97;
assign img[15755] = 97;
assign img[15756] = 97;
assign img[15757] = 97;
assign img[15758] = 105;
assign img[15759] = 96;
assign img[15760] = 97;
assign img[15761] = 112;
assign img[15762] = 107;
assign img[15763] = 104;
assign img[15764] = 105;
assign img[15765] = 105;
assign img[15766] = 105;
assign img[15767] = 128;
assign img[15768] = 106;
assign img[15769] = 109;
assign img[15770] = 106;
assign img[15771] = 100;
assign img[15772] = 109;
assign img[15773] = 104;
assign img[15774] = 105;
assign img[15775] = 99;
assign img[15776] = 108;
assign img[15777] = 128;
assign img[15778] = 101;
assign img[15779] = 128;
assign img[15780] = 108;
assign img[15781] = 112;
assign img[15782] = 128;
assign img[15783] = 109;
assign img[15784] = 128;
assign img[15785] = 105;
assign img[15786] = 102;
assign img[15787] = 128;
assign img[15788] = 105;
assign img[15789] = 105;
assign img[15790] = 105;
assign img[15791] = 128;
assign img[15792] = 111;
assign img[15793] = 108;
assign img[15794] = 104;
assign img[15795] = 104;
assign img[15796] = 105;
assign img[15797] = 105;
assign img[15798] = 112;
assign img[15799] = 102;
assign img[15800] = 108;
assign img[15801] = 112;
assign img[15802] = 104;
assign img[15803] = 128;
assign img[15804] = 103;
assign img[15805] = 106;
assign img[15806] = 128;
assign img[15807] = 110;
assign img[15808] = 104;
assign img[15809] = 109;
assign img[15810] = 104;
assign img[15811] = 105;
assign img[15812] = 114;
assign img[15813] = 108;
assign img[15814] = 108;
assign img[15815] = 109;
assign img[15816] = 108;
assign img[15817] = 110;
assign img[15818] = 108;
assign img[15819] = 104;
assign img[15820] = 100;
assign img[15821] = 96;
assign img[15822] = 100;
assign img[15823] = 90;
assign img[15824] = 90;
assign img[15825] = 88;
assign img[15826] = 86;
assign img[15827] = 96;
assign img[15828] = 90;
assign img[15829] = 88;
assign img[15830] = 88;
assign img[15831] = 88;
assign img[15832] = 79;
assign img[15833] = 81;
assign img[15834] = 92;
assign img[15835] = 84;
assign img[15836] = 84;
assign img[15837] = 88;
assign img[15838] = 87;
assign img[15839] = 87;
assign img[15840] = 85;
assign img[15841] = 88;
assign img[15842] = 92;
assign img[15843] = 88;
assign img[15844] = 82;
assign img[15845] = 83;
assign img[15846] = 86;
assign img[15847] = 86;
assign img[15848] = 82;
assign img[15849] = 87;
assign img[15850] = 88;
assign img[15851] = 96;
assign img[15852] = 81;
assign img[15853] = 88;
assign img[15854] = 82;
assign img[15855] = 82;
assign img[15856] = 93;
assign img[15857] = 80;
assign img[15858] = 81;
assign img[15859] = 83;
assign img[15860] = 76;
assign img[15861] = 80;
assign img[15862] = 80;
assign img[15863] = 84;
assign img[15864] = 84;
assign img[15865] = 78;
assign img[15866] = 84;
assign img[15867] = 73;
assign img[15868] = 79;
assign img[15869] = 79;
assign img[15870] = 83;
assign img[15871] = 84;
assign img[15872] = 82;
assign img[15873] = 96;
assign img[15874] = 90;
assign img[15875] = 91;
assign img[15876] = 91;
assign img[15877] = 100;
assign img[15878] = 102;
assign img[15879] = 96;
assign img[15880] = 97;
assign img[15881] = 100;
assign img[15882] = 96;
assign img[15883] = 100;
assign img[15884] = 98;
assign img[15885] = 98;
assign img[15886] = 96;
assign img[15887] = 99;
assign img[15888] = 97;
assign img[15889] = 104;
assign img[15890] = 104;
assign img[15891] = 128;
assign img[15892] = 128;
assign img[15893] = 128;
assign img[15894] = 113;
assign img[15895] = 113;
assign img[15896] = 107;
assign img[15897] = 128;
assign img[15898] = 105;
assign img[15899] = 113;
assign img[15900] = 104;
assign img[15901] = 128;
assign img[15902] = 128;
assign img[15903] = 112;
assign img[15904] = 128;
assign img[15905] = 112;
assign img[15906] = 128;
assign img[15907] = 128;
assign img[15908] = 105;
assign img[15909] = 113;
assign img[15910] = 128;
assign img[15911] = 109;
assign img[15912] = 112;
assign img[15913] = 128;
assign img[15914] = 109;
assign img[15915] = 128;
assign img[15916] = 128;
assign img[15917] = 109;
assign img[15918] = 128;
assign img[15919] = 105;
assign img[15920] = 128;
assign img[15921] = 112;
assign img[15922] = 128;
assign img[15923] = 105;
assign img[15924] = 105;
assign img[15925] = 111;
assign img[15926] = 128;
assign img[15927] = 128;
assign img[15928] = 109;
assign img[15929] = 110;
assign img[15930] = 111;
assign img[15931] = 128;
assign img[15932] = 128;
assign img[15933] = 110;
assign img[15934] = 108;
assign img[15935] = 128;
assign img[15936] = 109;
assign img[15937] = 128;
assign img[15938] = 128;
assign img[15939] = 128;
assign img[15940] = 113;
assign img[15941] = 107;
assign img[15942] = 105;
assign img[15943] = 112;
assign img[15944] = 108;
assign img[15945] = 104;
assign img[15946] = 105;
assign img[15947] = 99;
assign img[15948] = 106;
assign img[15949] = 101;
assign img[15950] = 96;
assign img[15951] = 100;
assign img[15952] = 104;
assign img[15953] = 94;
assign img[15954] = 92;
assign img[15955] = 96;
assign img[15956] = 94;
assign img[15957] = 95;
assign img[15958] = 92;
assign img[15959] = 86;
assign img[15960] = 84;
assign img[15961] = 92;
assign img[15962] = 94;
assign img[15963] = 88;
assign img[15964] = 94;
assign img[15965] = 92;
assign img[15966] = 86;
assign img[15967] = 92;
assign img[15968] = 87;
assign img[15969] = 92;
assign img[15970] = 85;
assign img[15971] = 88;
assign img[15972] = 89;
assign img[15973] = 96;
assign img[15974] = 90;
assign img[15975] = 96;
assign img[15976] = 87;
assign img[15977] = 88;
assign img[15978] = 85;
assign img[15979] = 87;
assign img[15980] = 92;
assign img[15981] = 88;
assign img[15982] = 90;
assign img[15983] = 96;
assign img[15984] = 86;
assign img[15985] = 84;
assign img[15986] = 94;
assign img[15987] = 88;
assign img[15988] = 92;
assign img[15989] = 84;
assign img[15990] = 86;
assign img[15991] = 87;
assign img[15992] = 86;
assign img[15993] = 84;
assign img[15994] = 79;
assign img[15995] = 79;
assign img[15996] = 86;
assign img[15997] = 96;
assign img[15998] = 92;
assign img[15999] = 87;
assign img[16000] = 84;
assign img[16001] = 109;
assign img[16002] = 96;
assign img[16003] = 102;
assign img[16004] = 96;
assign img[16005] = 96;
assign img[16006] = 96;
assign img[16007] = 102;
assign img[16008] = 98;
assign img[16009] = 112;
assign img[16010] = 105;
assign img[16011] = 103;
assign img[16012] = 96;
assign img[16013] = 128;
assign img[16014] = 101;
assign img[16015] = 110;
assign img[16016] = 108;
assign img[16017] = 128;
assign img[16018] = 128;
assign img[16019] = 113;
assign img[16020] = 111;
assign img[16021] = 128;
assign img[16022] = 128;
assign img[16023] = 128;
assign img[16024] = 128;
assign img[16025] = 128;
assign img[16026] = 128;
assign img[16027] = 129;
assign img[16028] = 129;
assign img[16029] = 128;
assign img[16030] = 129;
assign img[16031] = 128;
assign img[16032] = 128;
assign img[16033] = 128;
assign img[16034] = 128;
assign img[16035] = 128;
assign img[16036] = 129;
assign img[16037] = 128;
assign img[16038] = 128;
assign img[16039] = 128;
assign img[16040] = 128;
assign img[16041] = 128;
assign img[16042] = 128;
assign img[16043] = 128;
assign img[16044] = 128;
assign img[16045] = 128;
assign img[16046] = 128;
assign img[16047] = 128;
assign img[16048] = 128;
assign img[16049] = 128;
assign img[16050] = 129;
assign img[16051] = 128;
assign img[16052] = 128;
assign img[16053] = 128;
assign img[16054] = 128;
assign img[16055] = 128;
assign img[16056] = 128;
assign img[16057] = 133;
assign img[16058] = 128;
assign img[16059] = 129;
assign img[16060] = 129;
assign img[16061] = 128;
assign img[16062] = 128;
assign img[16063] = 129;
assign img[16064] = 128;
assign img[16065] = 129;
assign img[16066] = 128;
assign img[16067] = 129;
assign img[16068] = 128;
assign img[16069] = 128;
assign img[16070] = 128;
assign img[16071] = 113;
assign img[16072] = 100;
assign img[16073] = 105;
assign img[16074] = 100;
assign img[16075] = 104;
assign img[16076] = 97;
assign img[16077] = 98;
assign img[16078] = 100;
assign img[16079] = 104;
assign img[16080] = 98;
assign img[16081] = 108;
assign img[16082] = 96;
assign img[16083] = 102;
assign img[16084] = 100;
assign img[16085] = 96;
assign img[16086] = 103;
assign img[16087] = 94;
assign img[16088] = 98;
assign img[16089] = 102;
assign img[16090] = 102;
assign img[16091] = 98;
assign img[16092] = 98;
assign img[16093] = 96;
assign img[16094] = 98;
assign img[16095] = 96;
assign img[16096] = 96;
assign img[16097] = 96;
assign img[16098] = 100;
assign img[16099] = 96;
assign img[16100] = 96;
assign img[16101] = 96;
assign img[16102] = 96;
assign img[16103] = 92;
assign img[16104] = 96;
assign img[16105] = 97;
assign img[16106] = 96;
assign img[16107] = 97;
assign img[16108] = 93;
assign img[16109] = 95;
assign img[16110] = 97;
assign img[16111] = 97;
assign img[16112] = 96;
assign img[16113] = 96;
assign img[16114] = 91;
assign img[16115] = 92;
assign img[16116] = 96;
assign img[16117] = 96;
assign img[16118] = 90;
assign img[16119] = 87;
assign img[16120] = 102;
assign img[16121] = 96;
assign img[16122] = 87;
assign img[16123] = 90;
assign img[16124] = 98;
assign img[16125] = 97;
assign img[16126] = 98;
assign img[16127] = 96;
assign img[16128] = 87;
assign img[16129] = 104;
assign img[16130] = 128;
assign img[16131] = 112;
assign img[16132] = 112;
assign img[16133] = 128;
assign img[16134] = 110;
assign img[16135] = 128;
assign img[16136] = 111;
assign img[16137] = 116;
assign img[16138] = 112;
assign img[16139] = 128;
assign img[16140] = 115;
assign img[16141] = 109;
assign img[16142] = 105;
assign img[16143] = 128;
assign img[16144] = 109;
assign img[16145] = 113;
assign img[16146] = 128;
assign img[16147] = 128;
assign img[16148] = 128;
assign img[16149] = 129;
assign img[16150] = 113;
assign img[16151] = 128;
assign img[16152] = 128;
assign img[16153] = 113;
assign img[16154] = 128;
assign img[16155] = 128;
assign img[16156] = 128;
assign img[16157] = 128;
assign img[16158] = 128;
assign img[16159] = 128;
assign img[16160] = 128;
assign img[16161] = 129;
assign img[16162] = 129;
assign img[16163] = 128;
assign img[16164] = 128;
assign img[16165] = 128;
assign img[16166] = 129;
assign img[16167] = 131;
assign img[16168] = 129;
assign img[16169] = 129;
assign img[16170] = 138;
assign img[16171] = 129;
assign img[16172] = 129;
assign img[16173] = 128;
assign img[16174] = 130;
assign img[16175] = 130;
assign img[16176] = 128;
assign img[16177] = 128;
assign img[16178] = 128;
assign img[16179] = 128;
assign img[16180] = 128;
assign img[16181] = 128;
assign img[16182] = 128;
assign img[16183] = 128;
assign img[16184] = 128;
assign img[16185] = 128;
assign img[16186] = 129;
assign img[16187] = 128;
assign img[16188] = 128;
assign img[16189] = 129;
assign img[16190] = 129;
assign img[16191] = 128;
assign img[16192] = 128;
assign img[16193] = 128;
assign img[16194] = 128;
assign img[16195] = 112;
assign img[16196] = 128;
assign img[16197] = 128;
assign img[16198] = 111;
assign img[16199] = 128;
assign img[16200] = 128;
assign img[16201] = 128;
assign img[16202] = 109;
assign img[16203] = 110;
assign img[16204] = 128;
assign img[16205] = 97;
assign img[16206] = 107;
assign img[16207] = 108;
assign img[16208] = 105;
assign img[16209] = 111;
assign img[16210] = 100;
assign img[16211] = 128;
assign img[16212] = 105;
assign img[16213] = 100;
assign img[16214] = 104;
assign img[16215] = 108;
assign img[16216] = 108;
assign img[16217] = 128;
assign img[16218] = 108;
assign img[16219] = 112;
assign img[16220] = 110;
assign img[16221] = 111;
assign img[16222] = 108;
assign img[16223] = 100;
assign img[16224] = 108;
assign img[16225] = 128;
assign img[16226] = 128;
assign img[16227] = 110;
assign img[16228] = 108;
assign img[16229] = 112;
assign img[16230] = 108;
assign img[16231] = 96;
assign img[16232] = 104;
assign img[16233] = 109;
assign img[16234] = 100;
assign img[16235] = 103;
assign img[16236] = 108;
assign img[16237] = 101;
assign img[16238] = 108;
assign img[16239] = 109;
assign img[16240] = 100;
assign img[16241] = 108;
assign img[16242] = 100;
assign img[16243] = 104;
assign img[16244] = 100;
assign img[16245] = 104;
assign img[16246] = 108;
assign img[16247] = 104;
assign img[16248] = 99;
assign img[16249] = 100;
assign img[16250] = 108;
assign img[16251] = 102;
assign img[16252] = 100;
assign img[16253] = 100;
assign img[16254] = 108;
assign img[16255] = 108;
assign img[16256] = 98;
assign img[16257] = 128;
assign img[16258] = 128;
assign img[16259] = 128;
assign img[16260] = 129;
assign img[16261] = 128;
assign img[16262] = 128;
assign img[16263] = 128;
assign img[16264] = 128;
assign img[16265] = 129;
assign img[16266] = 128;
assign img[16267] = 128;
assign img[16268] = 129;
assign img[16269] = 128;
assign img[16270] = 128;
assign img[16271] = 129;
assign img[16272] = 128;
assign img[16273] = 129;
assign img[16274] = 128;
assign img[16275] = 128;
assign img[16276] = 128;
assign img[16277] = 128;
assign img[16278] = 129;
assign img[16279] = 128;
assign img[16280] = 128;
assign img[16281] = 128;
assign img[16282] = 128;
assign img[16283] = 128;
assign img[16284] = 128;
assign img[16285] = 128;
assign img[16286] = 128;
assign img[16287] = 129;
assign img[16288] = 128;
assign img[16289] = 136;
assign img[16290] = 128;
assign img[16291] = 128;
assign img[16292] = 129;
assign img[16293] = 128;
assign img[16294] = 129;
assign img[16295] = 128;
assign img[16296] = 129;
assign img[16297] = 129;
assign img[16298] = 128;
assign img[16299] = 131;
assign img[16300] = 132;
assign img[16301] = 129;
assign img[16302] = 128;
assign img[16303] = 128;
assign img[16304] = 129;
assign img[16305] = 129;
assign img[16306] = 128;
assign img[16307] = 129;
assign img[16308] = 129;
assign img[16309] = 128;
assign img[16310] = 128;
assign img[16311] = 128;
assign img[16312] = 129;
assign img[16313] = 129;
assign img[16314] = 128;
assign img[16315] = 128;
assign img[16316] = 128;
assign img[16317] = 128;
assign img[16318] = 131;
assign img[16319] = 132;
assign img[16320] = 129;
assign img[16321] = 129;
assign img[16322] = 128;
assign img[16323] = 128;
assign img[16324] = 128;
assign img[16325] = 128;
assign img[16326] = 128;
assign img[16327] = 128;
assign img[16328] = 128;
assign img[16329] = 128;
assign img[16330] = 128;
assign img[16331] = 128;
assign img[16332] = 128;
assign img[16333] = 128;
assign img[16334] = 128;
assign img[16335] = 128;
assign img[16336] = 128;
assign img[16337] = 128;
assign img[16338] = 128;
assign img[16339] = 128;
assign img[16340] = 128;
assign img[16341] = 128;
assign img[16342] = 129;
assign img[16343] = 128;
assign img[16344] = 128;
assign img[16345] = 128;
assign img[16346] = 128;
assign img[16347] = 128;
assign img[16348] = 128;
assign img[16349] = 128;
assign img[16350] = 128;
assign img[16351] = 128;
assign img[16352] = 128;
assign img[16353] = 128;
assign img[16354] = 128;
assign img[16355] = 128;
assign img[16356] = 128;
assign img[16357] = 128;
assign img[16358] = 128;
assign img[16359] = 128;
assign img[16360] = 128;
assign img[16361] = 128;
assign img[16362] = 129;
assign img[16363] = 128;
assign img[16364] = 128;
assign img[16365] = 128;
assign img[16366] = 128;
assign img[16367] = 128;
assign img[16368] = 128;
assign img[16369] = 128;
assign img[16370] = 128;
assign img[16371] = 128;
assign img[16372] = 128;
assign img[16373] = 112;
assign img[16374] = 128;
assign img[16375] = 128;
assign img[16376] = 128;
assign img[16377] = 128;
assign img[16378] = 128;
assign img[16379] = 128;
assign img[16380] = 128;
assign img[16381] = 128;
assign img[16382] = 129;
assign img[16383] = 128;

endmodule