// File:    fdct_tb.sv
// Author:  Lei Kuang
// Date:    17th June 2020
// @ Imperial College London

module fdct_tb;

logic        clk;
logic        nrst;
logic [7:0]  din;
logic        din_valid;
logic [7:0]  dout;
logic        dout_valid;

fdct dut(.*);

initial begin
    clk = '0;
    forever #5ns clk = ~clk;
end

logic [13:0] din_cnt;
logic [7:0]  img [16383:0];

initial begin
    nrst      = '0;
    din_cnt   = '0;
    din_valid = '0;
    
    @(posedge clk)
        nrst <= '1;
    
    forever begin
        @(posedge clk) begin
            din_valid <= ~din_valid;

            if(din_valid)
                din_cnt <= din_cnt + 1;
        end
    end
end

assign din = img[din_cnt];

initial begin
    byte temp;
    integer cnt = 0;
    
    forever @ (negedge clk) begin
        if(dout_valid) begin
            if(cnt % 64 == 0)
                 $write("MCU: %d\n", cnt >> 6);

            temp = dout;
            $write("%6d", temp);

            cnt = cnt + 1;
            if(cnt % 8 == 0)
                $write("\n");

        end
    end
end

// Debug
logic [5:0] pix_cnt;
logic [7:0] mcu_cnt;

logic end_of_mcu;
logic end_of_img;

assign end_of_mcu = pix_cnt=='1;
assign end_of_img = mcu_cnt=='1;

always_ff @ (posedge clk, negedge nrst)
    if(~nrst) begin
        pix_cnt <= '0;
        mcu_cnt <= '0;
    end
    else begin
        if(dout_valid)
            pix_cnt <= pix_cnt + 6'd1;
        if(end_of_mcu)
            mcu_cnt <= mcu_cnt + 8'd1; 
    end
    
assign img[    0] = 64;
assign img[    1] = 220;
assign img[    2] = 253;
assign img[    3] = 255;
assign img[    4] = 255;
assign img[    5] = 255;
assign img[    6] = 206;
assign img[    7] = 238;
assign img[    8] = 222;
assign img[    9] = 255;
assign img[   10] = 255;
assign img[   11] = 223;
assign img[   12] = 221;
assign img[   13] = 253;
assign img[   14] = 255;
assign img[   15] = 255;
assign img[   16] = 255;
assign img[   17] = 255;
assign img[   18] = 255;
assign img[   19] = 255;
assign img[   20] = 170;
assign img[   21] = 238;
assign img[   22] = 254;
assign img[   23] = 255;
assign img[   24] = 255;
assign img[   25] = 255;
assign img[   26] = 221;
assign img[   27] = 253;
assign img[   28] = 223;
assign img[   29] = 253;
assign img[   30] = 239;
assign img[   31] = 191;
assign img[   32] = 171;
assign img[   33] = 238;
assign img[   34] = 254;
assign img[   35] = 255;
assign img[   36] = 255;
assign img[   37] = 255;
assign img[   38] = 255;
assign img[   39] = 255;
assign img[   40] = 238;
assign img[   41] = 254;
assign img[   42] = 238;
assign img[   43] = 255;
assign img[   44] = 255;
assign img[   45] = 223;
assign img[   46] = 252;
assign img[   47] = 223;
assign img[   48] = 253;
assign img[   49] = 255;
assign img[   50] = 255;
assign img[   51] = 255;
assign img[   52] = 255;
assign img[   53] = 255;
assign img[   54] = 255;
assign img[   55] = 255;
assign img[   56] = 239;
assign img[   57] = 255;
assign img[   58] = 255;
assign img[   59] = 239;
assign img[   60] = 238;
assign img[   61] = 238;
assign img[   62] = 238;
assign img[   63] = 255;
assign img[   64] = 255;
assign img[   65] = 255;
assign img[   66] = 223;
assign img[   67] = 255;
assign img[   68] = 255;
assign img[   69] = 255;
assign img[   70] = 255;
assign img[   71] = 255;
assign img[   72] = 238;
assign img[   73] = 238;
assign img[   74] = 255;
assign img[   75] = 239;
assign img[   76] = 238;
assign img[   77] = 255;
assign img[   78] = 221;
assign img[   79] = 255;
assign img[   80] = 255;
assign img[   81] = 255;
assign img[   82] = 223;
assign img[   83] = 221;
assign img[   84] = 236;
assign img[   85] = 255;
assign img[   86] = 255;
assign img[   87] = 255;
assign img[   88] = 239;
assign img[   89] = 238;
assign img[   90] = 238;
assign img[   91] = 238;
assign img[   92] = 254;
assign img[   93] = 255;
assign img[   94] = 255;
assign img[   95] = 255;
assign img[   96] = 170;
assign img[   97] = 251;
assign img[   98] = 255;
assign img[   99] = 239;
assign img[  100] = 238;
assign img[  101] = 238;
assign img[  102] = 254;
assign img[  103] = 255;
assign img[  104] = 255;
assign img[  105] = 255;
assign img[  106] = 255;
assign img[  107] = 255;
assign img[  108] = 206;
assign img[  109] = 238;
assign img[  110] = 238;
assign img[  111] = 238;
assign img[  112] = 254;
assign img[  113] = 255;
assign img[  114] = 255;
assign img[  115] = 223;
assign img[  116] = 221;
assign img[  117] = 253;
assign img[  118] = 255;
assign img[  119] = 255;
assign img[  120] = 255;
assign img[  121] = 255;
assign img[  122] = 255;
assign img[  123] = 255;
assign img[  124] = 255;
assign img[  125] = 255;
assign img[  126] = 254;
assign img[  127] = 255;
assign img[  128] = 96;
assign img[  129] = 239;
assign img[  130] = 238;
assign img[  131] = 255;
assign img[  132] = 221;
assign img[  133] = 255;
assign img[  134] = 255;
assign img[  135] = 255;
assign img[  136] = 255;
assign img[  137] = 255;
assign img[  138] = 255;
assign img[  139] = 223;
assign img[  140] = 204;
assign img[  141] = 238;
assign img[  142] = 238;
assign img[  143] = 223;
assign img[  144] = 221;
assign img[  145] = 255;
assign img[  146] = 255;
assign img[  147] = 255;
assign img[  148] = 238;
assign img[  149] = 238;
assign img[  150] = 255;
assign img[  151] = 255;
assign img[  152] = 255;
assign img[  153] = 255;
assign img[  154] = 170;
assign img[  155] = 254;
assign img[  156] = 255;
assign img[  157] = 255;
assign img[  158] = 239;
assign img[  159] = 239;
assign img[  160] = 156;
assign img[  161] = 255;
assign img[  162] = 255;
assign img[  163] = 255;
assign img[  164] = 255;
assign img[  165] = 255;
assign img[  166] = 255;
assign img[  167] = 223;
assign img[  168] = 253;
assign img[  169] = 255;
assign img[  170] = 239;
assign img[  171] = 255;
assign img[  172] = 255;
assign img[  173] = 239;
assign img[  174] = 238;
assign img[  175] = 238;
assign img[  176] = 254;
assign img[  177] = 255;
assign img[  178] = 255;
assign img[  179] = 255;
assign img[  180] = 255;
assign img[  181] = 255;
assign img[  182] = 255;
assign img[  183] = 255;
assign img[  184] = 255;
assign img[  185] = 255;
assign img[  186] = 255;
assign img[  187] = 255;
assign img[  188] = 255;
assign img[  189] = 255;
assign img[  190] = 255;
assign img[  191] = 255;
assign img[  192] = 255;
assign img[  193] = 255;
assign img[  194] = 255;
assign img[  195] = 255;
assign img[  196] = 255;
assign img[  197] = 239;
assign img[  198] = 238;
assign img[  199] = 238;
assign img[  200] = 238;
assign img[  201] = 238;
assign img[  202] = 255;
assign img[  203] = 255;
assign img[  204] = 255;
assign img[  205] = 255;
assign img[  206] = 255;
assign img[  207] = 255;
assign img[  208] = 255;
assign img[  209] = 255;
assign img[  210] = 255;
assign img[  211] = 255;
assign img[  212] = 255;
assign img[  213] = 223;
assign img[  214] = 238;
assign img[  215] = 238;
assign img[  216] = 255;
assign img[  217] = 255;
assign img[  218] = 223;
assign img[  219] = 255;
assign img[  220] = 238;
assign img[  221] = 238;
assign img[  222] = 238;
assign img[  223] = 174;
assign img[  224] = 206;
assign img[  225] = 204;
assign img[  226] = 252;
assign img[  227] = 255;
assign img[  228] = 255;
assign img[  229] = 223;
assign img[  230] = 236;
assign img[  231] = 254;
assign img[  232] = 255;
assign img[  233] = 255;
assign img[  234] = 238;
assign img[  235] = 238;
assign img[  236] = 206;
assign img[  237] = 238;
assign img[  238] = 238;
assign img[  239] = 255;
assign img[  240] = 255;
assign img[  241] = 255;
assign img[  242] = 255;
assign img[  243] = 255;
assign img[  244] = 255;
assign img[  245] = 255;
assign img[  246] = 255;
assign img[  247] = 255;
assign img[  248] = 255;
assign img[  249] = 239;
assign img[  250] = 238;
assign img[  251] = 255;
assign img[  252] = 255;
assign img[  253] = 255;
assign img[  254] = 239;
assign img[  255] = 238;
assign img[  256] = 96;
assign img[  257] = 238;
assign img[  258] = 238;
assign img[  259] = 255;
assign img[  260] = 255;
assign img[  261] = 255;
assign img[  262] = 239;
assign img[  263] = 255;
assign img[  264] = 255;
assign img[  265] = 255;
assign img[  266] = 255;
assign img[  267] = 255;
assign img[  268] = 238;
assign img[  269] = 238;
assign img[  270] = 238;
assign img[  271] = 238;
assign img[  272] = 204;
assign img[  273] = 238;
assign img[  274] = 254;
assign img[  275] = 255;
assign img[  276] = 239;
assign img[  277] = 238;
assign img[  278] = 238;
assign img[  279] = 238;
assign img[  280] = 238;
assign img[  281] = 191;
assign img[  282] = 171;
assign img[  283] = 238;
assign img[  284] = 238;
assign img[  285] = 238;
assign img[  286] = 222;
assign img[  287] = 239;
assign img[  288] = 238;
assign img[  289] = 238;
assign img[  290] = 238;
assign img[  291] = 238;
assign img[  292] = 254;
assign img[  293] = 223;
assign img[  294] = 253;
assign img[  295] = 255;
assign img[  296] = 255;
assign img[  297] = 255;
assign img[  298] = 255;
assign img[  299] = 239;
assign img[  300] = 238;
assign img[  301] = 238;
assign img[  302] = 238;
assign img[  303] = 238;
assign img[  304] = 254;
assign img[  305] = 255;
assign img[  306] = 255;
assign img[  307] = 255;
assign img[  308] = 238;
assign img[  309] = 255;
assign img[  310] = 255;
assign img[  311] = 255;
assign img[  312] = 238;
assign img[  313] = 255;
assign img[  314] = 238;
assign img[  315] = 238;
assign img[  316] = 238;
assign img[  317] = 238;
assign img[  318] = 238;
assign img[  319] = 255;
assign img[  320] = 255;
assign img[  321] = 255;
assign img[  322] = 255;
assign img[  323] = 255;
assign img[  324] = 239;
assign img[  325] = 255;
assign img[  326] = 171;
assign img[  327] = 238;
assign img[  328] = 238;
assign img[  329] = 238;
assign img[  330] = 254;
assign img[  331] = 255;
assign img[  332] = 255;
assign img[  333] = 255;
assign img[  334] = 255;
assign img[  335] = 255;
assign img[  336] = 255;
assign img[  337] = 255;
assign img[  338] = 255;
assign img[  339] = 255;
assign img[  340] = 207;
assign img[  341] = 238;
assign img[  342] = 238;
assign img[  343] = 238;
assign img[  344] = 238;
assign img[  345] = 254;
assign img[  346] = 206;
assign img[  347] = 223;
assign img[  348] = 238;
assign img[  349] = 255;
assign img[  350] = 254;
assign img[  351] = 255;
assign img[  352] = 255;
assign img[  353] = 206;
assign img[  354] = 236;
assign img[  355] = 238;
assign img[  356] = 238;
assign img[  357] = 255;
assign img[  358] = 238;
assign img[  359] = 238;
assign img[  360] = 238;
assign img[  361] = 255;
assign img[  362] = 255;
assign img[  363] = 239;
assign img[  364] = 238;
assign img[  365] = 238;
assign img[  366] = 238;
assign img[  367] = 255;
assign img[  368] = 255;
assign img[  369] = 255;
assign img[  370] = 255;
assign img[  371] = 255;
assign img[  372] = 238;
assign img[  373] = 238;
assign img[  374] = 238;
assign img[  375] = 238;
assign img[  376] = 206;
assign img[  377] = 255;
assign img[  378] = 238;
assign img[  379] = 238;
assign img[  380] = 170;
assign img[  381] = 234;
assign img[  382] = 238;
assign img[  383] = 254;
assign img[  384] = 96;
assign img[  385] = 255;
assign img[  386] = 255;
assign img[  387] = 255;
assign img[  388] = 255;
assign img[  389] = 239;
assign img[  390] = 254;
assign img[  391] = 239;
assign img[  392] = 238;
assign img[  393] = 238;
assign img[  394] = 238;
assign img[  395] = 206;
assign img[  396] = 220;
assign img[  397] = 253;
assign img[  398] = 255;
assign img[  399] = 239;
assign img[  400] = 204;
assign img[  401] = 221;
assign img[  402] = 253;
assign img[  403] = 255;
assign img[  404] = 187;
assign img[  405] = 255;
assign img[  406] = 223;
assign img[  407] = 255;
assign img[  408] = 255;
assign img[  409] = 255;
assign img[  410] = 239;
assign img[  411] = 238;
assign img[  412] = 238;
assign img[  413] = 255;
assign img[  414] = 255;
assign img[  415] = 239;
assign img[  416] = 126;
assign img[  417] = 255;
assign img[  418] = 255;
assign img[  419] = 255;
assign img[  420] = 255;
assign img[  421] = 255;
assign img[  422] = 255;
assign img[  423] = 255;
assign img[  424] = 255;
assign img[  425] = 255;
assign img[  426] = 255;
assign img[  427] = 239;
assign img[  428] = 238;
assign img[  429] = 238;
assign img[  430] = 238;
assign img[  431] = 255;
assign img[  432] = 255;
assign img[  433] = 255;
assign img[  434] = 255;
assign img[  435] = 255;
assign img[  436] = 221;
assign img[  437] = 255;
assign img[  438] = 207;
assign img[  439] = 238;
assign img[  440] = 238;
assign img[  441] = 206;
assign img[  442] = 204;
assign img[  443] = 221;
assign img[  444] = 253;
assign img[  445] = 239;
assign img[  446] = 238;
assign img[  447] = 238;
assign img[  448] = 238;
assign img[  449] = 238;
assign img[  450] = 238;
assign img[  451] = 238;
assign img[  452] = 206;
assign img[  453] = 223;
assign img[  454] = 221;
assign img[  455] = 253;
assign img[  456] = 255;
assign img[  457] = 223;
assign img[  458] = 204;
assign img[  459] = 255;
assign img[  460] = 238;
assign img[  461] = 238;
assign img[  462] = 238;
assign img[  463] = 255;
assign img[  464] = 255;
assign img[  465] = 255;
assign img[  466] = 255;
assign img[  467] = 255;
assign img[  468] = 255;
assign img[  469] = 239;
assign img[  470] = 238;
assign img[  471] = 238;
assign img[  472] = 254;
assign img[  473] = 255;
assign img[  474] = 255;
assign img[  475] = 191;
assign img[  476] = 255;
assign img[  477] = 255;
assign img[  478] = 255;
assign img[  479] = 255;
assign img[  480] = 221;
assign img[  481] = 205;
assign img[  482] = 254;
assign img[  483] = 255;
assign img[  484] = 255;
assign img[  485] = 223;
assign img[  486] = 236;
assign img[  487] = 238;
assign img[  488] = 238;
assign img[  489] = 255;
assign img[  490] = 254;
assign img[  491] = 255;
assign img[  492] = 255;
assign img[  493] = 255;
assign img[  494] = 255;
assign img[  495] = 255;
assign img[  496] = 255;
assign img[  497] = 255;
assign img[  498] = 255;
assign img[  499] = 255;
assign img[  500] = 221;
assign img[  501] = 253;
assign img[  502] = 255;
assign img[  503] = 255;
assign img[  504] = 255;
assign img[  505] = 255;
assign img[  506] = 171;
assign img[  507] = 170;
assign img[  508] = 136;
assign img[  509] = 238;
assign img[  510] = 238;
assign img[  511] = 238;
assign img[  512] = 96;
assign img[  513] = 238;
assign img[  514] = 254;
assign img[  515] = 255;
assign img[  516] = 223;
assign img[  517] = 239;
assign img[  518] = 238;
assign img[  519] = 238;
assign img[  520] = 238;
assign img[  521] = 238;
assign img[  522] = 238;
assign img[  523] = 206;
assign img[  524] = 220;
assign img[  525] = 254;
assign img[  526] = 254;
assign img[  527] = 255;
assign img[  528] = 204;
assign img[  529] = 253;
assign img[  530] = 238;
assign img[  531] = 223;
assign img[  532] = 221;
assign img[  533] = 255;
assign img[  534] = 255;
assign img[  535] = 255;
assign img[  536] = 255;
assign img[  537] = 255;
assign img[  538] = 255;
assign img[  539] = 255;
assign img[  540] = 255;
assign img[  541] = 255;
assign img[  542] = 254;
assign img[  543] = 255;
assign img[  544] = 204;
assign img[  545] = 204;
assign img[  546] = 236;
assign img[  547] = 255;
assign img[  548] = 255;
assign img[  549] = 239;
assign img[  550] = 206;
assign img[  551] = 255;
assign img[  552] = 255;
assign img[  553] = 255;
assign img[  554] = 255;
assign img[  555] = 255;
assign img[  556] = 239;
assign img[  557] = 238;
assign img[  558] = 238;
assign img[  559] = 238;
assign img[  560] = 254;
assign img[  561] = 255;
assign img[  562] = 255;
assign img[  563] = 239;
assign img[  564] = 238;
assign img[  565] = 255;
assign img[  566] = 255;
assign img[  567] = 255;
assign img[  568] = 255;
assign img[  569] = 255;
assign img[  570] = 255;
assign img[  571] = 255;
assign img[  572] = 255;
assign img[  573] = 223;
assign img[  574] = 255;
assign img[  575] = 255;
assign img[  576] = 255;
assign img[  577] = 255;
assign img[  578] = 239;
assign img[  579] = 238;
assign img[  580] = 254;
assign img[  581] = 255;
assign img[  582] = 255;
assign img[  583] = 255;
assign img[  584] = 255;
assign img[  585] = 239;
assign img[  586] = 254;
assign img[  587] = 255;
assign img[  588] = 255;
assign img[  589] = 239;
assign img[  590] = 238;
assign img[  591] = 255;
assign img[  592] = 255;
assign img[  593] = 255;
assign img[  594] = 255;
assign img[  595] = 255;
assign img[  596] = 238;
assign img[  597] = 255;
assign img[  598] = 238;
assign img[  599] = 238;
assign img[  600] = 206;
assign img[  601] = 220;
assign img[  602] = 253;
assign img[  603] = 239;
assign img[  604] = 254;
assign img[  605] = 255;
assign img[  606] = 255;
assign img[  607] = 223;
assign img[  608] = 204;
assign img[  609] = 254;
assign img[  610] = 255;
assign img[  611] = 255;
assign img[  612] = 254;
assign img[  613] = 206;
assign img[  614] = 238;
assign img[  615] = 238;
assign img[  616] = 238;
assign img[  617] = 255;
assign img[  618] = 255;
assign img[  619] = 239;
assign img[  620] = 254;
assign img[  621] = 255;
assign img[  622] = 255;
assign img[  623] = 223;
assign img[  624] = 221;
assign img[  625] = 253;
assign img[  626] = 255;
assign img[  627] = 239;
assign img[  628] = 254;
assign img[  629] = 255;
assign img[  630] = 255;
assign img[  631] = 239;
assign img[  632] = 238;
assign img[  633] = 239;
assign img[  634] = 255;
assign img[  635] = 207;
assign img[  636] = 254;
assign img[  637] = 255;
assign img[  638] = 255;
assign img[  639] = 255;
assign img[  640] = 96;
assign img[  641] = 238;
assign img[  642] = 238;
assign img[  643] = 238;
assign img[  644] = 238;
assign img[  645] = 238;
assign img[  646] = 238;
assign img[  647] = 238;
assign img[  648] = 238;
assign img[  649] = 255;
assign img[  650] = 255;
assign img[  651] = 255;
assign img[  652] = 221;
assign img[  653] = 255;
assign img[  654] = 255;
assign img[  655] = 255;
assign img[  656] = 255;
assign img[  657] = 239;
assign img[  658] = 238;
assign img[  659] = 238;
assign img[  660] = 238;
assign img[  661] = 238;
assign img[  662] = 254;
assign img[  663] = 255;
assign img[  664] = 255;
assign img[  665] = 255;
assign img[  666] = 255;
assign img[  667] = 255;
assign img[  668] = 255;
assign img[  669] = 255;
assign img[  670] = 255;
assign img[  671] = 159;
assign img[  672] = 249;
assign img[  673] = 255;
assign img[  674] = 255;
assign img[  675] = 255;
assign img[  676] = 255;
assign img[  677] = 255;
assign img[  678] = 255;
assign img[  679] = 255;
assign img[  680] = 255;
assign img[  681] = 255;
assign img[  682] = 255;
assign img[  683] = 255;
assign img[  684] = 255;
assign img[  685] = 255;
assign img[  686] = 255;
assign img[  687] = 239;
assign img[  688] = 254;
assign img[  689] = 255;
assign img[  690] = 255;
assign img[  691] = 255;
assign img[  692] = 255;
assign img[  693] = 255;
assign img[  694] = 255;
assign img[  695] = 255;
assign img[  696] = 255;
assign img[  697] = 255;
assign img[  698] = 238;
assign img[  699] = 238;
assign img[  700] = 238;
assign img[  701] = 255;
assign img[  702] = 238;
assign img[  703] = 255;
assign img[  704] = 255;
assign img[  705] = 255;
assign img[  706] = 239;
assign img[  707] = 238;
assign img[  708] = 238;
assign img[  709] = 239;
assign img[  710] = 238;
assign img[  711] = 238;
assign img[  712] = 238;
assign img[  713] = 238;
assign img[  714] = 238;
assign img[  715] = 255;
assign img[  716] = 255;
assign img[  717] = 239;
assign img[  718] = 238;
assign img[  719] = 255;
assign img[  720] = 255;
assign img[  721] = 255;
assign img[  722] = 255;
assign img[  723] = 255;
assign img[  724] = 255;
assign img[  725] = 255;
assign img[  726] = 255;
assign img[  727] = 255;
assign img[  728] = 255;
assign img[  729] = 255;
assign img[  730] = 255;
assign img[  731] = 255;
assign img[  732] = 255;
assign img[  733] = 255;
assign img[  734] = 255;
assign img[  735] = 255;
assign img[  736] = 187;
assign img[  737] = 251;
assign img[  738] = 255;
assign img[  739] = 255;
assign img[  740] = 255;
assign img[  741] = 255;
assign img[  742] = 255;
assign img[  743] = 255;
assign img[  744] = 255;
assign img[  745] = 255;
assign img[  746] = 255;
assign img[  747] = 255;
assign img[  748] = 255;
assign img[  749] = 255;
assign img[  750] = 255;
assign img[  751] = 191;
assign img[  752] = 219;
assign img[  753] = 205;
assign img[  754] = 252;
assign img[  755] = 239;
assign img[  756] = 238;
assign img[  757] = 255;
assign img[  758] = 255;
assign img[  759] = 255;
assign img[  760] = 255;
assign img[  761] = 239;
assign img[  762] = 238;
assign img[  763] = 255;
assign img[  764] = 221;
assign img[  765] = 255;
assign img[  766] = 255;
assign img[  767] = 255;
assign img[  768] = 96;
assign img[  769] = 238;
assign img[  770] = 254;
assign img[  771] = 255;
assign img[  772] = 238;
assign img[  773] = 238;
assign img[  774] = 254;
assign img[  775] = 239;
assign img[  776] = 238;
assign img[  777] = 238;
assign img[  778] = 238;
assign img[  779] = 238;
assign img[  780] = 238;
assign img[  781] = 238;
assign img[  782] = 174;
assign img[  783] = 171;
assign img[  784] = 170;
assign img[  785] = 238;
assign img[  786] = 238;
assign img[  787] = 223;
assign img[  788] = 238;
assign img[  789] = 238;
assign img[  790] = 238;
assign img[  791] = 238;
assign img[  792] = 238;
assign img[  793] = 254;
assign img[  794] = 238;
assign img[  795] = 238;
assign img[  796] = 238;
assign img[  797] = 255;
assign img[  798] = 255;
assign img[  799] = 207;
assign img[  800] = 238;
assign img[  801] = 238;
assign img[  802] = 238;
assign img[  803] = 238;
assign img[  804] = 238;
assign img[  805] = 238;
assign img[  806] = 255;
assign img[  807] = 255;
assign img[  808] = 255;
assign img[  809] = 255;
assign img[  810] = 223;
assign img[  811] = 255;
assign img[  812] = 255;
assign img[  813] = 255;
assign img[  814] = 255;
assign img[  815] = 223;
assign img[  816] = 255;
assign img[  817] = 255;
assign img[  818] = 255;
assign img[  819] = 239;
assign img[  820] = 238;
assign img[  821] = 238;
assign img[  822] = 238;
assign img[  823] = 255;
assign img[  824] = 255;
assign img[  825] = 255;
assign img[  826] = 239;
assign img[  827] = 254;
assign img[  828] = 255;
assign img[  829] = 223;
assign img[  830] = 220;
assign img[  831] = 253;
assign img[  832] = 255;
assign img[  833] = 255;
assign img[  834] = 221;
assign img[  835] = 253;
assign img[  836] = 255;
assign img[  837] = 255;
assign img[  838] = 238;
assign img[  839] = 254;
assign img[  840] = 254;
assign img[  841] = 255;
assign img[  842] = 255;
assign img[  843] = 255;
assign img[  844] = 255;
assign img[  845] = 255;
assign img[  846] = 255;
assign img[  847] = 255;
assign img[  848] = 223;
assign img[  849] = 255;
assign img[  850] = 255;
assign img[  851] = 255;
assign img[  852] = 239;
assign img[  853] = 254;
assign img[  854] = 255;
assign img[  855] = 255;
assign img[  856] = 255;
assign img[  857] = 255;
assign img[  858] = 255;
assign img[  859] = 255;
assign img[  860] = 255;
assign img[  861] = 255;
assign img[  862] = 255;
assign img[  863] = 255;
assign img[  864] = 255;
assign img[  865] = 255;
assign img[  866] = 255;
assign img[  867] = 255;
assign img[  868] = 255;
assign img[  869] = 255;
assign img[  870] = 223;
assign img[  871] = 255;
assign img[  872] = 255;
assign img[  873] = 255;
assign img[  874] = 255;
assign img[  875] = 255;
assign img[  876] = 239;
assign img[  877] = 238;
assign img[  878] = 190;
assign img[  879] = 187;
assign img[  880] = 187;
assign img[  881] = 187;
assign img[  882] = 251;
assign img[  883] = 255;
assign img[  884] = 255;
assign img[  885] = 255;
assign img[  886] = 255;
assign img[  887] = 255;
assign img[  888] = 255;
assign img[  889] = 255;
assign img[  890] = 255;
assign img[  891] = 255;
assign img[  892] = 238;
assign img[  893] = 254;
assign img[  894] = 255;
assign img[  895] = 255;
assign img[  896] = 64;
assign img[  897] = 220;
assign img[  898] = 253;
assign img[  899] = 207;
assign img[  900] = 204;
assign img[  901] = 204;
assign img[  902] = 204;
assign img[  903] = 236;
assign img[  904] = 238;
assign img[  905] = 238;
assign img[  906] = 223;
assign img[  907] = 205;
assign img[  908] = 220;
assign img[  909] = 221;
assign img[  910] = 205;
assign img[  911] = 238;
assign img[  912] = 238;
assign img[  913] = 239;
assign img[  914] = 238;
assign img[  915] = 238;
assign img[  916] = 238;
assign img[  917] = 238;
assign img[  918] = 238;
assign img[  919] = 254;
assign img[  920] = 255;
assign img[  921] = 238;
assign img[  922] = 238;
assign img[  923] = 238;
assign img[  924] = 238;
assign img[  925] = 255;
assign img[  926] = 255;
assign img[  927] = 239;
assign img[  928] = 204;
assign img[  929] = 252;
assign img[  930] = 206;
assign img[  931] = 255;
assign img[  932] = 255;
assign img[  933] = 255;
assign img[  934] = 255;
assign img[  935] = 239;
assign img[  936] = 238;
assign img[  937] = 238;
assign img[  938] = 238;
assign img[  939] = 238;
assign img[  940] = 238;
assign img[  941] = 238;
assign img[  942] = 238;
assign img[  943] = 239;
assign img[  944] = 238;
assign img[  945] = 238;
assign img[  946] = 254;
assign img[  947] = 239;
assign img[  948] = 238;
assign img[  949] = 255;
assign img[  950] = 255;
assign img[  951] = 255;
assign img[  952] = 255;
assign img[  953] = 255;
assign img[  954] = 255;
assign img[  955] = 255;
assign img[  956] = 238;
assign img[  957] = 238;
assign img[  958] = 238;
assign img[  959] = 255;
assign img[  960] = 255;
assign img[  961] = 255;
assign img[  962] = 239;
assign img[  963] = 238;
assign img[  964] = 238;
assign img[  965] = 255;
assign img[  966] = 255;
assign img[  967] = 239;
assign img[  968] = 254;
assign img[  969] = 255;
assign img[  970] = 255;
assign img[  971] = 255;
assign img[  972] = 255;
assign img[  973] = 255;
assign img[  974] = 255;
assign img[  975] = 255;
assign img[  976] = 239;
assign img[  977] = 238;
assign img[  978] = 238;
assign img[  979] = 238;
assign img[  980] = 238;
assign img[  981] = 238;
assign img[  982] = 238;
assign img[  983] = 238;
assign img[  984] = 238;
assign img[  985] = 254;
assign img[  986] = 239;
assign img[  987] = 238;
assign img[  988] = 254;
assign img[  989] = 255;
assign img[  990] = 255;
assign img[  991] = 255;
assign img[  992] = 223;
assign img[  993] = 255;
assign img[  994] = 255;
assign img[  995] = 255;
assign img[  996] = 255;
assign img[  997] = 223;
assign img[  998] = 205;
assign img[  999] = 236;
assign img[ 1000] = 254;
assign img[ 1001] = 255;
assign img[ 1002] = 238;
assign img[ 1003] = 238;
assign img[ 1004] = 238;
assign img[ 1005] = 238;
assign img[ 1006] = 238;
assign img[ 1007] = 255;
assign img[ 1008] = 255;
assign img[ 1009] = 255;
assign img[ 1010] = 255;
assign img[ 1011] = 255;
assign img[ 1012] = 255;
assign img[ 1013] = 223;
assign img[ 1014] = 253;
assign img[ 1015] = 255;
assign img[ 1016] = 255;
assign img[ 1017] = 255;
assign img[ 1018] = 255;
assign img[ 1019] = 255;
assign img[ 1020] = 221;
assign img[ 1021] = 253;
assign img[ 1022] = 255;
assign img[ 1023] = 205;
assign img[ 1024] = 96;
assign img[ 1025] = 238;
assign img[ 1026] = 238;
assign img[ 1027] = 255;
assign img[ 1028] = 255;
assign img[ 1029] = 255;
assign img[ 1030] = 205;
assign img[ 1031] = 238;
assign img[ 1032] = 238;
assign img[ 1033] = 206;
assign img[ 1034] = 204;
assign img[ 1035] = 220;
assign img[ 1036] = 221;
assign img[ 1037] = 221;
assign img[ 1038] = 221;
assign img[ 1039] = 221;
assign img[ 1040] = 253;
assign img[ 1041] = 255;
assign img[ 1042] = 255;
assign img[ 1043] = 223;
assign img[ 1044] = 253;
assign img[ 1045] = 255;
assign img[ 1046] = 239;
assign img[ 1047] = 238;
assign img[ 1048] = 238;
assign img[ 1049] = 255;
assign img[ 1050] = 170;
assign img[ 1051] = 234;
assign img[ 1052] = 238;
assign img[ 1053] = 255;
assign img[ 1054] = 255;
assign img[ 1055] = 207;
assign img[ 1056] = 220;
assign img[ 1057] = 255;
assign img[ 1058] = 191;
assign img[ 1059] = 255;
assign img[ 1060] = 255;
assign img[ 1061] = 255;
assign img[ 1062] = 255;
assign img[ 1063] = 255;
assign img[ 1064] = 255;
assign img[ 1065] = 255;
assign img[ 1066] = 191;
assign img[ 1067] = 255;
assign img[ 1068] = 238;
assign img[ 1069] = 238;
assign img[ 1070] = 254;
assign img[ 1071] = 238;
assign img[ 1072] = 238;
assign img[ 1073] = 238;
assign img[ 1074] = 238;
assign img[ 1075] = 255;
assign img[ 1076] = 255;
assign img[ 1077] = 255;
assign img[ 1078] = 255;
assign img[ 1079] = 255;
assign img[ 1080] = 223;
assign img[ 1081] = 205;
assign img[ 1082] = 236;
assign img[ 1083] = 254;
assign img[ 1084] = 255;
assign img[ 1085] = 239;
assign img[ 1086] = 255;
assign img[ 1087] = 255;
assign img[ 1088] = 255;
assign img[ 1089] = 255;
assign img[ 1090] = 255;
assign img[ 1091] = 255;
assign img[ 1092] = 255;
assign img[ 1093] = 255;
assign img[ 1094] = 238;
assign img[ 1095] = 238;
assign img[ 1096] = 238;
assign img[ 1097] = 255;
assign img[ 1098] = 255;
assign img[ 1099] = 255;
assign img[ 1100] = 255;
assign img[ 1101] = 255;
assign img[ 1102] = 255;
assign img[ 1103] = 255;
assign img[ 1104] = 255;
assign img[ 1105] = 255;
assign img[ 1106] = 223;
assign img[ 1107] = 255;
assign img[ 1108] = 239;
assign img[ 1109] = 238;
assign img[ 1110] = 238;
assign img[ 1111] = 255;
assign img[ 1112] = 255;
assign img[ 1113] = 255;
assign img[ 1114] = 255;
assign img[ 1115] = 239;
assign img[ 1116] = 254;
assign img[ 1117] = 255;
assign img[ 1118] = 255;
assign img[ 1119] = 255;
assign img[ 1120] = 255;
assign img[ 1121] = 239;
assign img[ 1122] = 254;
assign img[ 1123] = 255;
assign img[ 1124] = 255;
assign img[ 1125] = 255;
assign img[ 1126] = 221;
assign img[ 1127] = 255;
assign img[ 1128] = 255;
assign img[ 1129] = 255;
assign img[ 1130] = 238;
assign img[ 1131] = 238;
assign img[ 1132] = 206;
assign img[ 1133] = 238;
assign img[ 1134] = 238;
assign img[ 1135] = 238;
assign img[ 1136] = 254;
assign img[ 1137] = 255;
assign img[ 1138] = 239;
assign img[ 1139] = 222;
assign img[ 1140] = 221;
assign img[ 1141] = 205;
assign img[ 1142] = 204;
assign img[ 1143] = 236;
assign img[ 1144] = 254;
assign img[ 1145] = 255;
assign img[ 1146] = 238;
assign img[ 1147] = 255;
assign img[ 1148] = 238;
assign img[ 1149] = 238;
assign img[ 1150] = 238;
assign img[ 1151] = 238;
assign img[ 1152] = 96;
assign img[ 1153] = 191;
assign img[ 1154] = 234;
assign img[ 1155] = 206;
assign img[ 1156] = 220;
assign img[ 1157] = 255;
assign img[ 1158] = 255;
assign img[ 1159] = 255;
assign img[ 1160] = 255;
assign img[ 1161] = 255;
assign img[ 1162] = 255;
assign img[ 1163] = 255;
assign img[ 1164] = 221;
assign img[ 1165] = 255;
assign img[ 1166] = 255;
assign img[ 1167] = 239;
assign img[ 1168] = 254;
assign img[ 1169] = 255;
assign img[ 1170] = 255;
assign img[ 1171] = 239;
assign img[ 1172] = 238;
assign img[ 1173] = 238;
assign img[ 1174] = 206;
assign img[ 1175] = 255;
assign img[ 1176] = 255;
assign img[ 1177] = 207;
assign img[ 1178] = 204;
assign img[ 1179] = 238;
assign img[ 1180] = 254;
assign img[ 1181] = 255;
assign img[ 1182] = 255;
assign img[ 1183] = 191;
assign img[ 1184] = 251;
assign img[ 1185] = 255;
assign img[ 1186] = 255;
assign img[ 1187] = 255;
assign img[ 1188] = 255;
assign img[ 1189] = 239;
assign img[ 1190] = 238;
assign img[ 1191] = 255;
assign img[ 1192] = 255;
assign img[ 1193] = 255;
assign img[ 1194] = 239;
assign img[ 1195] = 254;
assign img[ 1196] = 239;
assign img[ 1197] = 206;
assign img[ 1198] = 236;
assign img[ 1199] = 238;
assign img[ 1200] = 238;
assign img[ 1201] = 238;
assign img[ 1202] = 238;
assign img[ 1203] = 206;
assign img[ 1204] = 204;
assign img[ 1205] = 204;
assign img[ 1206] = 236;
assign img[ 1207] = 255;
assign img[ 1208] = 255;
assign img[ 1209] = 223;
assign img[ 1210] = 236;
assign img[ 1211] = 238;
assign img[ 1212] = 204;
assign img[ 1213] = 205;
assign img[ 1214] = 236;
assign img[ 1215] = 255;
assign img[ 1216] = 255;
assign img[ 1217] = 255;
assign img[ 1218] = 239;
assign img[ 1219] = 255;
assign img[ 1220] = 223;
assign img[ 1221] = 221;
assign img[ 1222] = 204;
assign img[ 1223] = 236;
assign img[ 1224] = 238;
assign img[ 1225] = 238;
assign img[ 1226] = 238;
assign img[ 1227] = 207;
assign img[ 1228] = 204;
assign img[ 1229] = 236;
assign img[ 1230] = 238;
assign img[ 1231] = 238;
assign img[ 1232] = 254;
assign img[ 1233] = 255;
assign img[ 1234] = 223;
assign img[ 1235] = 255;
assign img[ 1236] = 238;
assign img[ 1237] = 238;
assign img[ 1238] = 238;
assign img[ 1239] = 238;
assign img[ 1240] = 206;
assign img[ 1241] = 238;
assign img[ 1242] = 238;
assign img[ 1243] = 255;
assign img[ 1244] = 238;
assign img[ 1245] = 238;
assign img[ 1246] = 238;
assign img[ 1247] = 206;
assign img[ 1248] = 140;
assign img[ 1249] = 153;
assign img[ 1250] = 251;
assign img[ 1251] = 255;
assign img[ 1252] = 255;
assign img[ 1253] = 239;
assign img[ 1254] = 206;
assign img[ 1255] = 254;
assign img[ 1256] = 255;
assign img[ 1257] = 255;
assign img[ 1258] = 255;
assign img[ 1259] = 255;
assign img[ 1260] = 206;
assign img[ 1261] = 238;
assign img[ 1262] = 238;
assign img[ 1263] = 238;
assign img[ 1264] = 170;
assign img[ 1265] = 238;
assign img[ 1266] = 238;
assign img[ 1267] = 238;
assign img[ 1268] = 222;
assign img[ 1269] = 221;
assign img[ 1270] = 221;
assign img[ 1271] = 255;
assign img[ 1272] = 255;
assign img[ 1273] = 255;
assign img[ 1274] = 239;
assign img[ 1275] = 238;
assign img[ 1276] = 238;
assign img[ 1277] = 238;
assign img[ 1278] = 174;
assign img[ 1279] = 238;
assign img[ 1280] = 96;
assign img[ 1281] = 223;
assign img[ 1282] = 253;
assign img[ 1283] = 255;
assign img[ 1284] = 255;
assign img[ 1285] = 239;
assign img[ 1286] = 254;
assign img[ 1287] = 255;
assign img[ 1288] = 255;
assign img[ 1289] = 239;
assign img[ 1290] = 238;
assign img[ 1291] = 238;
assign img[ 1292] = 206;
assign img[ 1293] = 204;
assign img[ 1294] = 204;
assign img[ 1295] = 204;
assign img[ 1296] = 204;
assign img[ 1297] = 204;
assign img[ 1298] = 236;
assign img[ 1299] = 238;
assign img[ 1300] = 238;
assign img[ 1301] = 254;
assign img[ 1302] = 255;
assign img[ 1303] = 255;
assign img[ 1304] = 255;
assign img[ 1305] = 238;
assign img[ 1306] = 254;
assign img[ 1307] = 255;
assign img[ 1308] = 255;
assign img[ 1309] = 255;
assign img[ 1310] = 239;
assign img[ 1311] = 207;
assign img[ 1312] = 153;
assign img[ 1313] = 251;
assign img[ 1314] = 255;
assign img[ 1315] = 255;
assign img[ 1316] = 255;
assign img[ 1317] = 255;
assign img[ 1318] = 255;
assign img[ 1319] = 255;
assign img[ 1320] = 255;
assign img[ 1321] = 255;
assign img[ 1322] = 255;
assign img[ 1323] = 255;
assign img[ 1324] = 255;
assign img[ 1325] = 255;
assign img[ 1326] = 255;
assign img[ 1327] = 223;
assign img[ 1328] = 253;
assign img[ 1329] = 255;
assign img[ 1330] = 239;
assign img[ 1331] = 206;
assign img[ 1332] = 204;
assign img[ 1333] = 255;
assign img[ 1334] = 223;
assign img[ 1335] = 253;
assign img[ 1336] = 238;
assign img[ 1337] = 238;
assign img[ 1338] = 238;
assign img[ 1339] = 254;
assign img[ 1340] = 255;
assign img[ 1341] = 255;
assign img[ 1342] = 255;
assign img[ 1343] = 255;
assign img[ 1344] = 255;
assign img[ 1345] = 255;
assign img[ 1346] = 255;
assign img[ 1347] = 255;
assign img[ 1348] = 255;
assign img[ 1349] = 255;
assign img[ 1350] = 255;
assign img[ 1351] = 254;
assign img[ 1352] = 238;
assign img[ 1353] = 223;
assign img[ 1354] = 253;
assign img[ 1355] = 255;
assign img[ 1356] = 223;
assign img[ 1357] = 255;
assign img[ 1358] = 238;
assign img[ 1359] = 255;
assign img[ 1360] = 207;
assign img[ 1361] = 238;
assign img[ 1362] = 254;
assign img[ 1363] = 255;
assign img[ 1364] = 255;
assign img[ 1365] = 239;
assign img[ 1366] = 238;
assign img[ 1367] = 238;
assign img[ 1368] = 238;
assign img[ 1369] = 238;
assign img[ 1370] = 254;
assign img[ 1371] = 255;
assign img[ 1372] = 255;
assign img[ 1373] = 239;
assign img[ 1374] = 238;
assign img[ 1375] = 174;
assign img[ 1376] = 238;
assign img[ 1377] = 254;
assign img[ 1378] = 255;
assign img[ 1379] = 255;
assign img[ 1380] = 255;
assign img[ 1381] = 255;
assign img[ 1382] = 255;
assign img[ 1383] = 255;
assign img[ 1384] = 255;
assign img[ 1385] = 239;
assign img[ 1386] = 238;
assign img[ 1387] = 238;
assign img[ 1388] = 238;
assign img[ 1389] = 238;
assign img[ 1390] = 222;
assign img[ 1391] = 221;
assign img[ 1392] = 221;
assign img[ 1393] = 221;
assign img[ 1394] = 221;
assign img[ 1395] = 205;
assign img[ 1396] = 204;
assign img[ 1397] = 254;
assign img[ 1398] = 255;
assign img[ 1399] = 255;
assign img[ 1400] = 254;
assign img[ 1401] = 191;
assign img[ 1402] = 186;
assign img[ 1403] = 238;
assign img[ 1404] = 254;
assign img[ 1405] = 255;
assign img[ 1406] = 255;
assign img[ 1407] = 255;
assign img[ 1408] = 96;
assign img[ 1409] = 206;
assign img[ 1410] = 252;
assign img[ 1411] = 223;
assign img[ 1412] = 157;
assign img[ 1413] = 221;
assign img[ 1414] = 205;
assign img[ 1415] = 236;
assign img[ 1416] = 238;
assign img[ 1417] = 254;
assign img[ 1418] = 239;
assign img[ 1419] = 206;
assign img[ 1420] = 236;
assign img[ 1421] = 238;
assign img[ 1422] = 238;
assign img[ 1423] = 238;
assign img[ 1424] = 238;
assign img[ 1425] = 223;
assign img[ 1426] = 253;
assign img[ 1427] = 255;
assign img[ 1428] = 238;
assign img[ 1429] = 238;
assign img[ 1430] = 254;
assign img[ 1431] = 255;
assign img[ 1432] = 255;
assign img[ 1433] = 255;
assign img[ 1434] = 255;
assign img[ 1435] = 255;
assign img[ 1436] = 255;
assign img[ 1437] = 255;
assign img[ 1438] = 255;
assign img[ 1439] = 223;
assign img[ 1440] = 253;
assign img[ 1441] = 255;
assign img[ 1442] = 255;
assign img[ 1443] = 255;
assign img[ 1444] = 255;
assign img[ 1445] = 239;
assign img[ 1446] = 238;
assign img[ 1447] = 238;
assign img[ 1448] = 238;
assign img[ 1449] = 238;
assign img[ 1450] = 238;
assign img[ 1451] = 254;
assign img[ 1452] = 221;
assign img[ 1453] = 221;
assign img[ 1454] = 255;
assign img[ 1455] = 255;
assign img[ 1456] = 255;
assign img[ 1457] = 255;
assign img[ 1458] = 255;
assign img[ 1459] = 255;
assign img[ 1460] = 255;
assign img[ 1461] = 255;
assign img[ 1462] = 255;
assign img[ 1463] = 239;
assign img[ 1464] = 238;
assign img[ 1465] = 238;
assign img[ 1466] = 206;
assign img[ 1467] = 238;
assign img[ 1468] = 238;
assign img[ 1469] = 255;
assign img[ 1470] = 255;
assign img[ 1471] = 255;
assign img[ 1472] = 255;
assign img[ 1473] = 255;
assign img[ 1474] = 239;
assign img[ 1475] = 238;
assign img[ 1476] = 254;
assign img[ 1477] = 255;
assign img[ 1478] = 255;
assign img[ 1479] = 255;
assign img[ 1480] = 255;
assign img[ 1481] = 255;
assign img[ 1482] = 255;
assign img[ 1483] = 239;
assign img[ 1484] = 238;
assign img[ 1485] = 254;
assign img[ 1486] = 255;
assign img[ 1487] = 255;
assign img[ 1488] = 239;
assign img[ 1489] = 238;
assign img[ 1490] = 254;
assign img[ 1491] = 255;
assign img[ 1492] = 255;
assign img[ 1493] = 255;
assign img[ 1494] = 238;
assign img[ 1495] = 238;
assign img[ 1496] = 254;
assign img[ 1497] = 255;
assign img[ 1498] = 239;
assign img[ 1499] = 238;
assign img[ 1500] = 238;
assign img[ 1501] = 238;
assign img[ 1502] = 254;
assign img[ 1503] = 175;
assign img[ 1504] = 202;
assign img[ 1505] = 204;
assign img[ 1506] = 238;
assign img[ 1507] = 238;
assign img[ 1508] = 238;
assign img[ 1509] = 255;
assign img[ 1510] = 255;
assign img[ 1511] = 255;
assign img[ 1512] = 255;
assign img[ 1513] = 239;
assign img[ 1514] = 238;
assign img[ 1515] = 239;
assign img[ 1516] = 238;
assign img[ 1517] = 254;
assign img[ 1518] = 255;
assign img[ 1519] = 255;
assign img[ 1520] = 255;
assign img[ 1521] = 239;
assign img[ 1522] = 238;
assign img[ 1523] = 238;
assign img[ 1524] = 206;
assign img[ 1525] = 206;
assign img[ 1526] = 255;
assign img[ 1527] = 255;
assign img[ 1528] = 238;
assign img[ 1529] = 255;
assign img[ 1530] = 221;
assign img[ 1531] = 221;
assign img[ 1532] = 253;
assign img[ 1533] = 255;
assign img[ 1534] = 207;
assign img[ 1535] = 236;
assign img[ 1536] = 112;
assign img[ 1537] = 239;
assign img[ 1538] = 238;
assign img[ 1539] = 239;
assign img[ 1540] = 255;
assign img[ 1541] = 255;
assign img[ 1542] = 255;
assign img[ 1543] = 255;
assign img[ 1544] = 255;
assign img[ 1545] = 255;
assign img[ 1546] = 255;
assign img[ 1547] = 255;
assign img[ 1548] = 255;
assign img[ 1549] = 255;
assign img[ 1550] = 255;
assign img[ 1551] = 255;
assign img[ 1552] = 255;
assign img[ 1553] = 255;
assign img[ 1554] = 255;
assign img[ 1555] = 255;
assign img[ 1556] = 187;
assign img[ 1557] = 255;
assign img[ 1558] = 239;
assign img[ 1559] = 238;
assign img[ 1560] = 238;
assign img[ 1561] = 239;
assign img[ 1562] = 238;
assign img[ 1563] = 238;
assign img[ 1564] = 238;
assign img[ 1565] = 255;
assign img[ 1566] = 239;
assign img[ 1567] = 206;
assign img[ 1568] = 252;
assign img[ 1569] = 255;
assign img[ 1570] = 207;
assign img[ 1571] = 238;
assign img[ 1572] = 238;
assign img[ 1573] = 222;
assign img[ 1574] = 221;
assign img[ 1575] = 255;
assign img[ 1576] = 255;
assign img[ 1577] = 255;
assign img[ 1578] = 255;
assign img[ 1579] = 255;
assign img[ 1580] = 239;
assign img[ 1581] = 255;
assign img[ 1582] = 255;
assign img[ 1583] = 239;
assign img[ 1584] = 238;
assign img[ 1585] = 238;
assign img[ 1586] = 238;
assign img[ 1587] = 238;
assign img[ 1588] = 238;
assign img[ 1589] = 254;
assign img[ 1590] = 255;
assign img[ 1591] = 255;
assign img[ 1592] = 255;
assign img[ 1593] = 255;
assign img[ 1594] = 239;
assign img[ 1595] = 238;
assign img[ 1596] = 238;
assign img[ 1597] = 238;
assign img[ 1598] = 238;
assign img[ 1599] = 255;
assign img[ 1600] = 255;
assign img[ 1601] = 255;
assign img[ 1602] = 255;
assign img[ 1603] = 255;
assign img[ 1604] = 255;
assign img[ 1605] = 255;
assign img[ 1606] = 221;
assign img[ 1607] = 255;
assign img[ 1608] = 221;
assign img[ 1609] = 255;
assign img[ 1610] = 255;
assign img[ 1611] = 239;
assign img[ 1612] = 238;
assign img[ 1613] = 254;
assign img[ 1614] = 255;
assign img[ 1615] = 255;
assign img[ 1616] = 223;
assign img[ 1617] = 255;
assign img[ 1618] = 255;
assign img[ 1619] = 255;
assign img[ 1620] = 238;
assign img[ 1621] = 238;
assign img[ 1622] = 238;
assign img[ 1623] = 238;
assign img[ 1624] = 254;
assign img[ 1625] = 255;
assign img[ 1626] = 221;
assign img[ 1627] = 253;
assign img[ 1628] = 238;
assign img[ 1629] = 206;
assign img[ 1630] = 254;
assign img[ 1631] = 191;
assign img[ 1632] = 255;
assign img[ 1633] = 255;
assign img[ 1634] = 255;
assign img[ 1635] = 255;
assign img[ 1636] = 255;
assign img[ 1637] = 255;
assign img[ 1638] = 239;
assign img[ 1639] = 238;
assign img[ 1640] = 238;
assign img[ 1641] = 239;
assign img[ 1642] = 238;
assign img[ 1643] = 238;
assign img[ 1644] = 254;
assign img[ 1645] = 255;
assign img[ 1646] = 255;
assign img[ 1647] = 255;
assign img[ 1648] = 255;
assign img[ 1649] = 255;
assign img[ 1650] = 255;
assign img[ 1651] = 255;
assign img[ 1652] = 239;
assign img[ 1653] = 238;
assign img[ 1654] = 238;
assign img[ 1655] = 238;
assign img[ 1656] = 238;
assign img[ 1657] = 238;
assign img[ 1658] = 238;
assign img[ 1659] = 255;
assign img[ 1660] = 205;
assign img[ 1661] = 238;
assign img[ 1662] = 238;
assign img[ 1663] = 254;
assign img[ 1664] = 96;
assign img[ 1665] = 223;
assign img[ 1666] = 253;
assign img[ 1667] = 255;
assign img[ 1668] = 221;
assign img[ 1669] = 221;
assign img[ 1670] = 221;
assign img[ 1671] = 221;
assign img[ 1672] = 253;
assign img[ 1673] = 255;
assign img[ 1674] = 255;
assign img[ 1675] = 239;
assign img[ 1676] = 238;
assign img[ 1677] = 238;
assign img[ 1678] = 238;
assign img[ 1679] = 238;
assign img[ 1680] = 204;
assign img[ 1681] = 238;
assign img[ 1682] = 238;
assign img[ 1683] = 255;
assign img[ 1684] = 255;
assign img[ 1685] = 255;
assign img[ 1686] = 255;
assign img[ 1687] = 255;
assign img[ 1688] = 255;
assign img[ 1689] = 239;
assign img[ 1690] = 238;
assign img[ 1691] = 238;
assign img[ 1692] = 238;
assign img[ 1693] = 255;
assign img[ 1694] = 255;
assign img[ 1695] = 255;
assign img[ 1696] = 255;
assign img[ 1697] = 223;
assign img[ 1698] = 236;
assign img[ 1699] = 255;
assign img[ 1700] = 239;
assign img[ 1701] = 238;
assign img[ 1702] = 238;
assign img[ 1703] = 255;
assign img[ 1704] = 255;
assign img[ 1705] = 255;
assign img[ 1706] = 255;
assign img[ 1707] = 255;
assign img[ 1708] = 255;
assign img[ 1709] = 255;
assign img[ 1710] = 255;
assign img[ 1711] = 223;
assign img[ 1712] = 253;
assign img[ 1713] = 255;
assign img[ 1714] = 255;
assign img[ 1715] = 255;
assign img[ 1716] = 223;
assign img[ 1717] = 221;
assign img[ 1718] = 253;
assign img[ 1719] = 255;
assign img[ 1720] = 239;
assign img[ 1721] = 255;
assign img[ 1722] = 239;
assign img[ 1723] = 238;
assign img[ 1724] = 238;
assign img[ 1725] = 238;
assign img[ 1726] = 238;
assign img[ 1727] = 255;
assign img[ 1728] = 255;
assign img[ 1729] = 255;
assign img[ 1730] = 255;
assign img[ 1731] = 255;
assign img[ 1732] = 255;
assign img[ 1733] = 255;
assign img[ 1734] = 204;
assign img[ 1735] = 221;
assign img[ 1736] = 253;
assign img[ 1737] = 255;
assign img[ 1738] = 255;
assign img[ 1739] = 255;
assign img[ 1740] = 255;
assign img[ 1741] = 255;
assign img[ 1742] = 255;
assign img[ 1743] = 255;
assign img[ 1744] = 223;
assign img[ 1745] = 255;
assign img[ 1746] = 255;
assign img[ 1747] = 255;
assign img[ 1748] = 255;
assign img[ 1749] = 255;
assign img[ 1750] = 255;
assign img[ 1751] = 255;
assign img[ 1752] = 223;
assign img[ 1753] = 255;
assign img[ 1754] = 191;
assign img[ 1755] = 187;
assign img[ 1756] = 234;
assign img[ 1757] = 238;
assign img[ 1758] = 238;
assign img[ 1759] = 254;
assign img[ 1760] = 187;
assign img[ 1761] = 251;
assign img[ 1762] = 238;
assign img[ 1763] = 255;
assign img[ 1764] = 238;
assign img[ 1765] = 255;
assign img[ 1766] = 223;
assign img[ 1767] = 255;
assign img[ 1768] = 238;
assign img[ 1769] = 255;
assign img[ 1770] = 238;
assign img[ 1771] = 255;
assign img[ 1772] = 238;
assign img[ 1773] = 255;
assign img[ 1774] = 254;
assign img[ 1775] = 255;
assign img[ 1776] = 255;
assign img[ 1777] = 255;
assign img[ 1778] = 255;
assign img[ 1779] = 239;
assign img[ 1780] = 254;
assign img[ 1781] = 255;
assign img[ 1782] = 254;
assign img[ 1783] = 255;
assign img[ 1784] = 255;
assign img[ 1785] = 175;
assign img[ 1786] = 187;
assign img[ 1787] = 207;
assign img[ 1788] = 204;
assign img[ 1789] = 236;
assign img[ 1790] = 238;
assign img[ 1791] = 238;
assign img[ 1792] = 96;
assign img[ 1793] = 206;
assign img[ 1794] = 252;
assign img[ 1795] = 255;
assign img[ 1796] = 223;
assign img[ 1797] = 253;
assign img[ 1798] = 255;
assign img[ 1799] = 255;
assign img[ 1800] = 255;
assign img[ 1801] = 255;
assign img[ 1802] = 239;
assign img[ 1803] = 238;
assign img[ 1804] = 238;
assign img[ 1805] = 238;
assign img[ 1806] = 238;
assign img[ 1807] = 207;
assign img[ 1808] = 236;
assign img[ 1809] = 238;
assign img[ 1810] = 238;
assign img[ 1811] = 223;
assign img[ 1812] = 238;
assign img[ 1813] = 238;
assign img[ 1814] = 254;
assign img[ 1815] = 255;
assign img[ 1816] = 255;
assign img[ 1817] = 255;
assign img[ 1818] = 187;
assign img[ 1819] = 255;
assign img[ 1820] = 238;
assign img[ 1821] = 255;
assign img[ 1822] = 254;
assign img[ 1823] = 238;
assign img[ 1824] = 238;
assign img[ 1825] = 238;
assign img[ 1826] = 238;
assign img[ 1827] = 238;
assign img[ 1828] = 238;
assign img[ 1829] = 254;
assign img[ 1830] = 255;
assign img[ 1831] = 239;
assign img[ 1832] = 238;
assign img[ 1833] = 238;
assign img[ 1834] = 238;
assign img[ 1835] = 238;
assign img[ 1836] = 238;
assign img[ 1837] = 239;
assign img[ 1838] = 238;
assign img[ 1839] = 255;
assign img[ 1840] = 255;
assign img[ 1841] = 255;
assign img[ 1842] = 255;
assign img[ 1843] = 239;
assign img[ 1844] = 238;
assign img[ 1845] = 255;
assign img[ 1846] = 255;
assign img[ 1847] = 255;
assign img[ 1848] = 255;
assign img[ 1849] = 255;
assign img[ 1850] = 255;
assign img[ 1851] = 255;
assign img[ 1852] = 255;
assign img[ 1853] = 255;
assign img[ 1854] = 255;
assign img[ 1855] = 255;
assign img[ 1856] = 255;
assign img[ 1857] = 255;
assign img[ 1858] = 255;
assign img[ 1859] = 255;
assign img[ 1860] = 255;
assign img[ 1861] = 239;
assign img[ 1862] = 238;
assign img[ 1863] = 255;
assign img[ 1864] = 255;
assign img[ 1865] = 255;
assign img[ 1866] = 255;
assign img[ 1867] = 255;
assign img[ 1868] = 223;
assign img[ 1869] = 255;
assign img[ 1870] = 255;
assign img[ 1871] = 255;
assign img[ 1872] = 255;
assign img[ 1873] = 255;
assign img[ 1874] = 239;
assign img[ 1875] = 223;
assign img[ 1876] = 221;
assign img[ 1877] = 255;
assign img[ 1878] = 255;
assign img[ 1879] = 255;
assign img[ 1880] = 239;
assign img[ 1881] = 238;
assign img[ 1882] = 238;
assign img[ 1883] = 238;
assign img[ 1884] = 238;
assign img[ 1885] = 238;
assign img[ 1886] = 238;
assign img[ 1887] = 255;
assign img[ 1888] = 221;
assign img[ 1889] = 237;
assign img[ 1890] = 238;
assign img[ 1891] = 238;
assign img[ 1892] = 238;
assign img[ 1893] = 238;
assign img[ 1894] = 254;
assign img[ 1895] = 255;
assign img[ 1896] = 255;
assign img[ 1897] = 239;
assign img[ 1898] = 238;
assign img[ 1899] = 238;
assign img[ 1900] = 206;
assign img[ 1901] = 238;
assign img[ 1902] = 254;
assign img[ 1903] = 255;
assign img[ 1904] = 255;
assign img[ 1905] = 255;
assign img[ 1906] = 255;
assign img[ 1907] = 255;
assign img[ 1908] = 238;
assign img[ 1909] = 238;
assign img[ 1910] = 238;
assign img[ 1911] = 238;
assign img[ 1912] = 238;
assign img[ 1913] = 238;
assign img[ 1914] = 238;
assign img[ 1915] = 206;
assign img[ 1916] = 220;
assign img[ 1917] = 255;
assign img[ 1918] = 223;
assign img[ 1919] = 253;
assign img[ 1920] = 96;
assign img[ 1921] = 238;
assign img[ 1922] = 238;
assign img[ 1923] = 238;
assign img[ 1924] = 206;
assign img[ 1925] = 204;
assign img[ 1926] = 252;
assign img[ 1927] = 255;
assign img[ 1928] = 255;
assign img[ 1929] = 255;
assign img[ 1930] = 255;
assign img[ 1931] = 191;
assign img[ 1932] = 251;
assign img[ 1933] = 255;
assign img[ 1934] = 223;
assign img[ 1935] = 223;
assign img[ 1936] = 255;
assign img[ 1937] = 237;
assign img[ 1938] = 238;
assign img[ 1939] = 238;
assign img[ 1940] = 204;
assign img[ 1941] = 238;
assign img[ 1942] = 238;
assign img[ 1943] = 238;
assign img[ 1944] = 238;
assign img[ 1945] = 223;
assign img[ 1946] = 221;
assign img[ 1947] = 221;
assign img[ 1948] = 204;
assign img[ 1949] = 254;
assign img[ 1950] = 206;
assign img[ 1951] = 252;
assign img[ 1952] = 255;
assign img[ 1953] = 255;
assign img[ 1954] = 255;
assign img[ 1955] = 255;
assign img[ 1956] = 223;
assign img[ 1957] = 221;
assign img[ 1958] = 253;
assign img[ 1959] = 207;
assign img[ 1960] = 236;
assign img[ 1961] = 255;
assign img[ 1962] = 221;
assign img[ 1963] = 253;
assign img[ 1964] = 238;
assign img[ 1965] = 206;
assign img[ 1966] = 236;
assign img[ 1967] = 255;
assign img[ 1968] = 255;
assign img[ 1969] = 255;
assign img[ 1970] = 239;
assign img[ 1971] = 238;
assign img[ 1972] = 206;
assign img[ 1973] = 238;
assign img[ 1974] = 206;
assign img[ 1975] = 238;
assign img[ 1976] = 238;
assign img[ 1977] = 255;
assign img[ 1978] = 255;
assign img[ 1979] = 255;
assign img[ 1980] = 255;
assign img[ 1981] = 255;
assign img[ 1982] = 255;
assign img[ 1983] = 255;
assign img[ 1984] = 255;
assign img[ 1985] = 255;
assign img[ 1986] = 255;
assign img[ 1987] = 255;
assign img[ 1988] = 255;
assign img[ 1989] = 255;
assign img[ 1990] = 255;
assign img[ 1991] = 255;
assign img[ 1992] = 255;
assign img[ 1993] = 239;
assign img[ 1994] = 238;
assign img[ 1995] = 239;
assign img[ 1996] = 255;
assign img[ 1997] = 255;
assign img[ 1998] = 238;
assign img[ 1999] = 255;
assign img[ 2000] = 255;
assign img[ 2001] = 255;
assign img[ 2002] = 223;
assign img[ 2003] = 221;
assign img[ 2004] = 237;
assign img[ 2005] = 206;
assign img[ 2006] = 204;
assign img[ 2007] = 238;
assign img[ 2008] = 238;
assign img[ 2009] = 255;
assign img[ 2010] = 255;
assign img[ 2011] = 207;
assign img[ 2012] = 252;
assign img[ 2013] = 255;
assign img[ 2014] = 255;
assign img[ 2015] = 255;
assign img[ 2016] = 255;
assign img[ 2017] = 255;
assign img[ 2018] = 255;
assign img[ 2019] = 239;
assign img[ 2020] = 238;
assign img[ 2021] = 238;
assign img[ 2022] = 204;
assign img[ 2023] = 236;
assign img[ 2024] = 254;
assign img[ 2025] = 255;
assign img[ 2026] = 255;
assign img[ 2027] = 239;
assign img[ 2028] = 238;
assign img[ 2029] = 238;
assign img[ 2030] = 238;
assign img[ 2031] = 238;
assign img[ 2032] = 238;
assign img[ 2033] = 238;
assign img[ 2034] = 220;
assign img[ 2035] = 255;
assign img[ 2036] = 157;
assign img[ 2037] = 137;
assign img[ 2038] = 232;
assign img[ 2039] = 238;
assign img[ 2040] = 238;
assign img[ 2041] = 238;
assign img[ 2042] = 238;
assign img[ 2043] = 255;
assign img[ 2044] = 221;
assign img[ 2045] = 255;
assign img[ 2046] = 255;
assign img[ 2047] = 255;
assign img[ 2048] = 96;
assign img[ 2049] = 207;
assign img[ 2050] = 253;
assign img[ 2051] = 255;
assign img[ 2052] = 255;
assign img[ 2053] = 255;
assign img[ 2054] = 191;
assign img[ 2055] = 254;
assign img[ 2056] = 254;
assign img[ 2057] = 255;
assign img[ 2058] = 238;
assign img[ 2059] = 238;
assign img[ 2060] = 206;
assign img[ 2061] = 204;
assign img[ 2062] = 204;
assign img[ 2063] = 204;
assign img[ 2064] = 204;
assign img[ 2065] = 204;
assign img[ 2066] = 236;
assign img[ 2067] = 191;
assign img[ 2068] = 155;
assign img[ 2069] = 255;
assign img[ 2070] = 239;
assign img[ 2071] = 255;
assign img[ 2072] = 255;
assign img[ 2073] = 255;
assign img[ 2074] = 187;
assign img[ 2075] = 255;
assign img[ 2076] = 255;
assign img[ 2077] = 255;
assign img[ 2078] = 255;
assign img[ 2079] = 255;
assign img[ 2080] = 103;
assign img[ 2081] = 230;
assign img[ 2082] = 238;
assign img[ 2083] = 255;
assign img[ 2084] = 223;
assign img[ 2085] = 255;
assign img[ 2086] = 238;
assign img[ 2087] = 238;
assign img[ 2088] = 238;
assign img[ 2089] = 238;
assign img[ 2090] = 190;
assign img[ 2091] = 171;
assign img[ 2092] = 170;
assign img[ 2093] = 238;
assign img[ 2094] = 238;
assign img[ 2095] = 238;
assign img[ 2096] = 238;
assign img[ 2097] = 238;
assign img[ 2098] = 238;
assign img[ 2099] = 255;
assign img[ 2100] = 255;
assign img[ 2101] = 255;
assign img[ 2102] = 255;
assign img[ 2103] = 239;
assign img[ 2104] = 238;
assign img[ 2105] = 238;
assign img[ 2106] = 238;
assign img[ 2107] = 238;
assign img[ 2108] = 238;
assign img[ 2109] = 255;
assign img[ 2110] = 255;
assign img[ 2111] = 255;
assign img[ 2112] = 255;
assign img[ 2113] = 255;
assign img[ 2114] = 191;
assign img[ 2115] = 255;
assign img[ 2116] = 255;
assign img[ 2117] = 255;
assign img[ 2118] = 238;
assign img[ 2119] = 238;
assign img[ 2120] = 254;
assign img[ 2121] = 255;
assign img[ 2122] = 254;
assign img[ 2123] = 255;
assign img[ 2124] = 255;
assign img[ 2125] = 255;
assign img[ 2126] = 255;
assign img[ 2127] = 255;
assign img[ 2128] = 255;
assign img[ 2129] = 255;
assign img[ 2130] = 255;
assign img[ 2131] = 255;
assign img[ 2132] = 238;
assign img[ 2133] = 174;
assign img[ 2134] = 234;
assign img[ 2135] = 238;
assign img[ 2136] = 238;
assign img[ 2137] = 238;
assign img[ 2138] = 238;
assign img[ 2139] = 206;
assign img[ 2140] = 252;
assign img[ 2141] = 255;
assign img[ 2142] = 255;
assign img[ 2143] = 255;
assign img[ 2144] = 187;
assign img[ 2145] = 119;
assign img[ 2146] = 247;
assign img[ 2147] = 255;
assign img[ 2148] = 255;
assign img[ 2149] = 239;
assign img[ 2150] = 254;
assign img[ 2151] = 255;
assign img[ 2152] = 255;
assign img[ 2153] = 255;
assign img[ 2154] = 238;
assign img[ 2155] = 255;
assign img[ 2156] = 221;
assign img[ 2157] = 255;
assign img[ 2158] = 255;
assign img[ 2159] = 255;
assign img[ 2160] = 223;
assign img[ 2161] = 221;
assign img[ 2162] = 221;
assign img[ 2163] = 221;
assign img[ 2164] = 237;
assign img[ 2165] = 255;
assign img[ 2166] = 221;
assign img[ 2167] = 255;
assign img[ 2168] = 255;
assign img[ 2169] = 239;
assign img[ 2170] = 255;
assign img[ 2171] = 255;
assign img[ 2172] = 255;
assign img[ 2173] = 255;
assign img[ 2174] = 239;
assign img[ 2175] = 238;
assign img[ 2176] = 96;
assign img[ 2177] = 238;
assign img[ 2178] = 238;
assign img[ 2179] = 238;
assign img[ 2180] = 254;
assign img[ 2181] = 255;
assign img[ 2182] = 207;
assign img[ 2183] = 238;
assign img[ 2184] = 238;
assign img[ 2185] = 238;
assign img[ 2186] = 238;
assign img[ 2187] = 238;
assign img[ 2188] = 222;
assign img[ 2189] = 255;
assign img[ 2190] = 159;
assign img[ 2191] = 205;
assign img[ 2192] = 236;
assign img[ 2193] = 206;
assign img[ 2194] = 236;
assign img[ 2195] = 174;
assign img[ 2196] = 170;
assign img[ 2197] = 238;
assign img[ 2198] = 238;
assign img[ 2199] = 255;
assign img[ 2200] = 255;
assign img[ 2201] = 255;
assign img[ 2202] = 255;
assign img[ 2203] = 255;
assign img[ 2204] = 255;
assign img[ 2205] = 255;
assign img[ 2206] = 255;
assign img[ 2207] = 191;
assign img[ 2208] = 187;
assign img[ 2209] = 251;
assign img[ 2210] = 255;
assign img[ 2211] = 223;
assign img[ 2212] = 255;
assign img[ 2213] = 255;
assign img[ 2214] = 255;
assign img[ 2215] = 255;
assign img[ 2216] = 255;
assign img[ 2217] = 255;
assign img[ 2218] = 239;
assign img[ 2219] = 238;
assign img[ 2220] = 238;
assign img[ 2221] = 238;
assign img[ 2222] = 238;
assign img[ 2223] = 238;
assign img[ 2224] = 254;
assign img[ 2225] = 239;
assign img[ 2226] = 238;
assign img[ 2227] = 238;
assign img[ 2228] = 204;
assign img[ 2229] = 238;
assign img[ 2230] = 238;
assign img[ 2231] = 238;
assign img[ 2232] = 238;
assign img[ 2233] = 239;
assign img[ 2234] = 238;
assign img[ 2235] = 238;
assign img[ 2236] = 238;
assign img[ 2237] = 255;
assign img[ 2238] = 255;
assign img[ 2239] = 255;
assign img[ 2240] = 255;
assign img[ 2241] = 255;
assign img[ 2242] = 255;
assign img[ 2243] = 254;
assign img[ 2244] = 238;
assign img[ 2245] = 255;
assign img[ 2246] = 239;
assign img[ 2247] = 238;
assign img[ 2248] = 238;
assign img[ 2249] = 238;
assign img[ 2250] = 238;
assign img[ 2251] = 255;
assign img[ 2252] = 238;
assign img[ 2253] = 254;
assign img[ 2254] = 255;
assign img[ 2255] = 255;
assign img[ 2256] = 255;
assign img[ 2257] = 255;
assign img[ 2258] = 255;
assign img[ 2259] = 239;
assign img[ 2260] = 238;
assign img[ 2261] = 175;
assign img[ 2262] = 238;
assign img[ 2263] = 238;
assign img[ 2264] = 238;
assign img[ 2265] = 238;
assign img[ 2266] = 238;
assign img[ 2267] = 238;
assign img[ 2268] = 206;
assign img[ 2269] = 238;
assign img[ 2270] = 238;
assign img[ 2271] = 174;
assign img[ 2272] = 170;
assign img[ 2273] = 187;
assign img[ 2274] = 251;
assign img[ 2275] = 239;
assign img[ 2276] = 238;
assign img[ 2277] = 238;
assign img[ 2278] = 238;
assign img[ 2279] = 238;
assign img[ 2280] = 254;
assign img[ 2281] = 255;
assign img[ 2282] = 255;
assign img[ 2283] = 255;
assign img[ 2284] = 255;
assign img[ 2285] = 255;
assign img[ 2286] = 255;
assign img[ 2287] = 255;
assign img[ 2288] = 223;
assign img[ 2289] = 223;
assign img[ 2290] = 239;
assign img[ 2291] = 223;
assign img[ 2292] = 157;
assign img[ 2293] = 221;
assign img[ 2294] = 221;
assign img[ 2295] = 255;
assign img[ 2296] = 255;
assign img[ 2297] = 223;
assign img[ 2298] = 204;
assign img[ 2299] = 221;
assign img[ 2300] = 253;
assign img[ 2301] = 255;
assign img[ 2302] = 255;
assign img[ 2303] = 255;
assign img[ 2304] = 96;
assign img[ 2305] = 238;
assign img[ 2306] = 238;
assign img[ 2307] = 238;
assign img[ 2308] = 250;
assign img[ 2309] = 255;
assign img[ 2310] = 223;
assign img[ 2311] = 255;
assign img[ 2312] = 255;
assign img[ 2313] = 255;
assign img[ 2314] = 238;
assign img[ 2315] = 222;
assign img[ 2316] = 253;
assign img[ 2317] = 254;
assign img[ 2318] = 239;
assign img[ 2319] = 206;
assign img[ 2320] = 220;
assign img[ 2321] = 253;
assign img[ 2322] = 238;
assign img[ 2323] = 255;
assign img[ 2324] = 255;
assign img[ 2325] = 255;
assign img[ 2326] = 255;
assign img[ 2327] = 255;
assign img[ 2328] = 239;
assign img[ 2329] = 255;
assign img[ 2330] = 187;
assign img[ 2331] = 255;
assign img[ 2332] = 238;
assign img[ 2333] = 255;
assign img[ 2334] = 255;
assign img[ 2335] = 207;
assign img[ 2336] = 204;
assign img[ 2337] = 238;
assign img[ 2338] = 238;
assign img[ 2339] = 255;
assign img[ 2340] = 223;
assign img[ 2341] = 205;
assign img[ 2342] = 204;
assign img[ 2343] = 204;
assign img[ 2344] = 252;
assign img[ 2345] = 255;
assign img[ 2346] = 255;
assign img[ 2347] = 255;
assign img[ 2348] = 255;
assign img[ 2349] = 238;
assign img[ 2350] = 238;
assign img[ 2351] = 239;
assign img[ 2352] = 255;
assign img[ 2353] = 255;
assign img[ 2354] = 239;
assign img[ 2355] = 254;
assign img[ 2356] = 255;
assign img[ 2357] = 255;
assign img[ 2358] = 255;
assign img[ 2359] = 255;
assign img[ 2360] = 255;
assign img[ 2361] = 255;
assign img[ 2362] = 239;
assign img[ 2363] = 255;
assign img[ 2364] = 255;
assign img[ 2365] = 255;
assign img[ 2366] = 255;
assign img[ 2367] = 255;
assign img[ 2368] = 255;
assign img[ 2369] = 255;
assign img[ 2370] = 223;
assign img[ 2371] = 255;
assign img[ 2372] = 255;
assign img[ 2373] = 239;
assign img[ 2374] = 238;
assign img[ 2375] = 238;
assign img[ 2376] = 238;
assign img[ 2377] = 238;
assign img[ 2378] = 255;
assign img[ 2379] = 255;
assign img[ 2380] = 255;
assign img[ 2381] = 255;
assign img[ 2382] = 255;
assign img[ 2383] = 255;
assign img[ 2384] = 255;
assign img[ 2385] = 255;
assign img[ 2386] = 255;
assign img[ 2387] = 223;
assign img[ 2388] = 253;
assign img[ 2389] = 223;
assign img[ 2390] = 253;
assign img[ 2391] = 255;
assign img[ 2392] = 255;
assign img[ 2393] = 223;
assign img[ 2394] = 221;
assign img[ 2395] = 221;
assign img[ 2396] = 253;
assign img[ 2397] = 255;
assign img[ 2398] = 255;
assign img[ 2399] = 255;
assign img[ 2400] = 255;
assign img[ 2401] = 239;
assign img[ 2402] = 254;
assign img[ 2403] = 255;
assign img[ 2404] = 239;
assign img[ 2405] = 238;
assign img[ 2406] = 238;
assign img[ 2407] = 206;
assign img[ 2408] = 236;
assign img[ 2409] = 238;
assign img[ 2410] = 238;
assign img[ 2411] = 238;
assign img[ 2412] = 206;
assign img[ 2413] = 238;
assign img[ 2414] = 238;
assign img[ 2415] = 238;
assign img[ 2416] = 238;
assign img[ 2417] = 238;
assign img[ 2418] = 238;
assign img[ 2419] = 238;
assign img[ 2420] = 238;
assign img[ 2421] = 255;
assign img[ 2422] = 238;
assign img[ 2423] = 238;
assign img[ 2424] = 238;
assign img[ 2425] = 238;
assign img[ 2426] = 238;
assign img[ 2427] = 238;
assign img[ 2428] = 254;
assign img[ 2429] = 255;
assign img[ 2430] = 255;
assign img[ 2431] = 255;
assign img[ 2432] = 96;
assign img[ 2433] = 206;
assign img[ 2434] = 252;
assign img[ 2435] = 239;
assign img[ 2436] = 220;
assign img[ 2437] = 253;
assign img[ 2438] = 207;
assign img[ 2439] = 204;
assign img[ 2440] = 236;
assign img[ 2441] = 238;
assign img[ 2442] = 254;
assign img[ 2443] = 255;
assign img[ 2444] = 221;
assign img[ 2445] = 221;
assign img[ 2446] = 255;
assign img[ 2447] = 223;
assign img[ 2448] = 221;
assign img[ 2449] = 255;
assign img[ 2450] = 255;
assign img[ 2451] = 255;
assign img[ 2452] = 221;
assign img[ 2453] = 255;
assign img[ 2454] = 255;
assign img[ 2455] = 255;
assign img[ 2456] = 238;
assign img[ 2457] = 223;
assign img[ 2458] = 253;
assign img[ 2459] = 255;
assign img[ 2460] = 255;
assign img[ 2461] = 255;
assign img[ 2462] = 255;
assign img[ 2463] = 175;
assign img[ 2464] = 138;
assign img[ 2465] = 255;
assign img[ 2466] = 255;
assign img[ 2467] = 255;
assign img[ 2468] = 223;
assign img[ 2469] = 221;
assign img[ 2470] = 253;
assign img[ 2471] = 207;
assign img[ 2472] = 236;
assign img[ 2473] = 238;
assign img[ 2474] = 238;
assign img[ 2475] = 191;
assign img[ 2476] = 239;
assign img[ 2477] = 238;
assign img[ 2478] = 238;
assign img[ 2479] = 238;
assign img[ 2480] = 238;
assign img[ 2481] = 238;
assign img[ 2482] = 254;
assign img[ 2483] = 255;
assign img[ 2484] = 221;
assign img[ 2485] = 253;
assign img[ 2486] = 255;
assign img[ 2487] = 255;
assign img[ 2488] = 255;
assign img[ 2489] = 191;
assign img[ 2490] = 187;
assign img[ 2491] = 187;
assign img[ 2492] = 250;
assign img[ 2493] = 223;
assign img[ 2494] = 255;
assign img[ 2495] = 255;
assign img[ 2496] = 255;
assign img[ 2497] = 255;
assign img[ 2498] = 255;
assign img[ 2499] = 255;
assign img[ 2500] = 255;
assign img[ 2501] = 255;
assign img[ 2502] = 191;
assign img[ 2503] = 187;
assign img[ 2504] = 251;
assign img[ 2505] = 255;
assign img[ 2506] = 255;
assign img[ 2507] = 207;
assign img[ 2508] = 204;
assign img[ 2509] = 236;
assign img[ 2510] = 238;
assign img[ 2511] = 238;
assign img[ 2512] = 238;
assign img[ 2513] = 254;
assign img[ 2514] = 255;
assign img[ 2515] = 238;
assign img[ 2516] = 204;
assign img[ 2517] = 255;
assign img[ 2518] = 255;
assign img[ 2519] = 255;
assign img[ 2520] = 255;
assign img[ 2521] = 255;
assign img[ 2522] = 255;
assign img[ 2523] = 207;
assign img[ 2524] = 238;
assign img[ 2525] = 238;
assign img[ 2526] = 254;
assign img[ 2527] = 239;
assign img[ 2528] = 254;
assign img[ 2529] = 239;
assign img[ 2530] = 254;
assign img[ 2531] = 255;
assign img[ 2532] = 255;
assign img[ 2533] = 255;
assign img[ 2534] = 239;
assign img[ 2535] = 238;
assign img[ 2536] = 238;
assign img[ 2537] = 238;
assign img[ 2538] = 238;
assign img[ 2539] = 239;
assign img[ 2540] = 238;
assign img[ 2541] = 238;
assign img[ 2542] = 238;
assign img[ 2543] = 238;
assign img[ 2544] = 254;
assign img[ 2545] = 255;
assign img[ 2546] = 255;
assign img[ 2547] = 255;
assign img[ 2548] = 255;
assign img[ 2549] = 255;
assign img[ 2550] = 255;
assign img[ 2551] = 255;
assign img[ 2552] = 255;
assign img[ 2553] = 207;
assign img[ 2554] = 238;
assign img[ 2555] = 206;
assign img[ 2556] = 204;
assign img[ 2557] = 253;
assign img[ 2558] = 255;
assign img[ 2559] = 255;
assign img[ 2560] = 96;
assign img[ 2561] = 206;
assign img[ 2562] = 236;
assign img[ 2563] = 238;
assign img[ 2564] = 238;
assign img[ 2565] = 238;
assign img[ 2566] = 254;
assign img[ 2567] = 255;
assign img[ 2568] = 255;
assign img[ 2569] = 255;
assign img[ 2570] = 255;
assign img[ 2571] = 255;
assign img[ 2572] = 255;
assign img[ 2573] = 255;
assign img[ 2574] = 255;
assign img[ 2575] = 207;
assign img[ 2576] = 204;
assign img[ 2577] = 238;
assign img[ 2578] = 238;
assign img[ 2579] = 255;
assign img[ 2580] = 187;
assign img[ 2581] = 251;
assign img[ 2582] = 207;
assign img[ 2583] = 238;
assign img[ 2584] = 238;
assign img[ 2585] = 239;
assign img[ 2586] = 238;
assign img[ 2587] = 238;
assign img[ 2588] = 238;
assign img[ 2589] = 238;
assign img[ 2590] = 254;
assign img[ 2591] = 206;
assign img[ 2592] = 204;
assign img[ 2593] = 254;
assign img[ 2594] = 255;
assign img[ 2595] = 255;
assign img[ 2596] = 238;
assign img[ 2597] = 255;
assign img[ 2598] = 238;
assign img[ 2599] = 255;
assign img[ 2600] = 238;
assign img[ 2601] = 255;
assign img[ 2602] = 254;
assign img[ 2603] = 255;
assign img[ 2604] = 238;
assign img[ 2605] = 239;
assign img[ 2606] = 238;
assign img[ 2607] = 255;
assign img[ 2608] = 255;
assign img[ 2609] = 255;
assign img[ 2610] = 255;
assign img[ 2611] = 255;
assign img[ 2612] = 255;
assign img[ 2613] = 255;
assign img[ 2614] = 255;
assign img[ 2615] = 255;
assign img[ 2616] = 255;
assign img[ 2617] = 255;
assign img[ 2618] = 239;
assign img[ 2619] = 238;
assign img[ 2620] = 238;
assign img[ 2621] = 222;
assign img[ 2622] = 253;
assign img[ 2623] = 255;
assign img[ 2624] = 255;
assign img[ 2625] = 255;
assign img[ 2626] = 223;
assign img[ 2627] = 221;
assign img[ 2628] = 236;
assign img[ 2629] = 255;
assign img[ 2630] = 238;
assign img[ 2631] = 238;
assign img[ 2632] = 238;
assign img[ 2633] = 238;
assign img[ 2634] = 238;
assign img[ 2635] = 238;
assign img[ 2636] = 238;
assign img[ 2637] = 238;
assign img[ 2638] = 238;
assign img[ 2639] = 255;
assign img[ 2640] = 239;
assign img[ 2641] = 238;
assign img[ 2642] = 238;
assign img[ 2643] = 238;
assign img[ 2644] = 238;
assign img[ 2645] = 238;
assign img[ 2646] = 238;
assign img[ 2647] = 238;
assign img[ 2648] = 254;
assign img[ 2649] = 255;
assign img[ 2650] = 255;
assign img[ 2651] = 255;
assign img[ 2652] = 255;
assign img[ 2653] = 255;
assign img[ 2654] = 255;
assign img[ 2655] = 255;
assign img[ 2656] = 255;
assign img[ 2657] = 239;
assign img[ 2658] = 238;
assign img[ 2659] = 238;
assign img[ 2660] = 238;
assign img[ 2661] = 238;
assign img[ 2662] = 238;
assign img[ 2663] = 238;
assign img[ 2664] = 238;
assign img[ 2665] = 239;
assign img[ 2666] = 238;
assign img[ 2667] = 238;
assign img[ 2668] = 138;
assign img[ 2669] = 238;
assign img[ 2670] = 238;
assign img[ 2671] = 238;
assign img[ 2672] = 238;
assign img[ 2673] = 238;
assign img[ 2674] = 254;
assign img[ 2675] = 255;
assign img[ 2676] = 171;
assign img[ 2677] = 238;
assign img[ 2678] = 238;
assign img[ 2679] = 238;
assign img[ 2680] = 238;
assign img[ 2681] = 206;
assign img[ 2682] = 220;
assign img[ 2683] = 221;
assign img[ 2684] = 221;
assign img[ 2685] = 255;
assign img[ 2686] = 223;
assign img[ 2687] = 253;
assign img[ 2688] = 96;
assign img[ 2689] = 238;
assign img[ 2690] = 238;
assign img[ 2691] = 255;
assign img[ 2692] = 221;
assign img[ 2693] = 255;
assign img[ 2694] = 223;
assign img[ 2695] = 255;
assign img[ 2696] = 255;
assign img[ 2697] = 255;
assign img[ 2698] = 255;
assign img[ 2699] = 223;
assign img[ 2700] = 221;
assign img[ 2701] = 255;
assign img[ 2702] = 239;
assign img[ 2703] = 238;
assign img[ 2704] = 220;
assign img[ 2705] = 221;
assign img[ 2706] = 236;
assign img[ 2707] = 223;
assign img[ 2708] = 236;
assign img[ 2709] = 238;
assign img[ 2710] = 238;
assign img[ 2711] = 238;
assign img[ 2712] = 254;
assign img[ 2713] = 255;
assign img[ 2714] = 170;
assign img[ 2715] = 238;
assign img[ 2716] = 254;
assign img[ 2717] = 255;
assign img[ 2718] = 255;
assign img[ 2719] = 255;
assign img[ 2720] = 255;
assign img[ 2721] = 255;
assign img[ 2722] = 255;
assign img[ 2723] = 255;
assign img[ 2724] = 255;
assign img[ 2725] = 255;
assign img[ 2726] = 239;
assign img[ 2727] = 238;
assign img[ 2728] = 238;
assign img[ 2729] = 238;
assign img[ 2730] = 238;
assign img[ 2731] = 254;
assign img[ 2732] = 255;
assign img[ 2733] = 207;
assign img[ 2734] = 236;
assign img[ 2735] = 238;
assign img[ 2736] = 254;
assign img[ 2737] = 255;
assign img[ 2738] = 255;
assign img[ 2739] = 255;
assign img[ 2740] = 239;
assign img[ 2741] = 238;
assign img[ 2742] = 238;
assign img[ 2743] = 238;
assign img[ 2744] = 238;
assign img[ 2745] = 238;
assign img[ 2746] = 238;
assign img[ 2747] = 255;
assign img[ 2748] = 238;
assign img[ 2749] = 238;
assign img[ 2750] = 238;
assign img[ 2751] = 255;
assign img[ 2752] = 255;
assign img[ 2753] = 255;
assign img[ 2754] = 239;
assign img[ 2755] = 238;
assign img[ 2756] = 238;
assign img[ 2757] = 238;
assign img[ 2758] = 238;
assign img[ 2759] = 238;
assign img[ 2760] = 255;
assign img[ 2761] = 255;
assign img[ 2762] = 255;
assign img[ 2763] = 255;
assign img[ 2764] = 238;
assign img[ 2765] = 238;
assign img[ 2766] = 238;
assign img[ 2767] = 255;
assign img[ 2768] = 255;
assign img[ 2769] = 255;
assign img[ 2770] = 255;
assign img[ 2771] = 255;
assign img[ 2772] = 255;
assign img[ 2773] = 255;
assign img[ 2774] = 238;
assign img[ 2775] = 238;
assign img[ 2776] = 206;
assign img[ 2777] = 204;
assign img[ 2778] = 236;
assign img[ 2779] = 238;
assign img[ 2780] = 238;
assign img[ 2781] = 238;
assign img[ 2782] = 238;
assign img[ 2783] = 190;
assign img[ 2784] = 187;
assign img[ 2785] = 235;
assign img[ 2786] = 254;
assign img[ 2787] = 255;
assign img[ 2788] = 255;
assign img[ 2789] = 255;
assign img[ 2790] = 238;
assign img[ 2791] = 238;
assign img[ 2792] = 238;
assign img[ 2793] = 238;
assign img[ 2794] = 238;
assign img[ 2795] = 238;
assign img[ 2796] = 206;
assign img[ 2797] = 238;
assign img[ 2798] = 238;
assign img[ 2799] = 238;
assign img[ 2800] = 238;
assign img[ 2801] = 238;
assign img[ 2802] = 238;
assign img[ 2803] = 255;
assign img[ 2804] = 255;
assign img[ 2805] = 255;
assign img[ 2806] = 255;
assign img[ 2807] = 255;
assign img[ 2808] = 255;
assign img[ 2809] = 239;
assign img[ 2810] = 238;
assign img[ 2811] = 255;
assign img[ 2812] = 255;
assign img[ 2813] = 255;
assign img[ 2814] = 255;
assign img[ 2815] = 255;
assign img[ 2816] = 0;
assign img[ 2817] = 136;
assign img[ 2818] = 232;
assign img[ 2819] = 238;
assign img[ 2820] = 238;
assign img[ 2821] = 238;
assign img[ 2822] = 238;
assign img[ 2823] = 238;
assign img[ 2824] = 238;
assign img[ 2825] = 238;
assign img[ 2826] = 238;
assign img[ 2827] = 223;
assign img[ 2828] = 255;
assign img[ 2829] = 238;
assign img[ 2830] = 238;
assign img[ 2831] = 223;
assign img[ 2832] = 221;
assign img[ 2833] = 253;
assign img[ 2834] = 253;
assign img[ 2835] = 255;
assign img[ 2836] = 221;
assign img[ 2837] = 239;
assign img[ 2838] = 238;
assign img[ 2839] = 239;
assign img[ 2840] = 238;
assign img[ 2841] = 238;
assign img[ 2842] = 238;
assign img[ 2843] = 238;
assign img[ 2844] = 238;
assign img[ 2845] = 255;
assign img[ 2846] = 223;
assign img[ 2847] = 221;
assign img[ 2848] = 221;
assign img[ 2849] = 255;
assign img[ 2850] = 255;
assign img[ 2851] = 255;
assign img[ 2852] = 239;
assign img[ 2853] = 254;
assign img[ 2854] = 255;
assign img[ 2855] = 238;
assign img[ 2856] = 204;
assign img[ 2857] = 236;
assign img[ 2858] = 238;
assign img[ 2859] = 238;
assign img[ 2860] = 238;
assign img[ 2861] = 255;
assign img[ 2862] = 255;
assign img[ 2863] = 255;
assign img[ 2864] = 255;
assign img[ 2865] = 255;
assign img[ 2866] = 191;
assign img[ 2867] = 187;
assign img[ 2868] = 251;
assign img[ 2869] = 255;
assign img[ 2870] = 207;
assign img[ 2871] = 238;
assign img[ 2872] = 238;
assign img[ 2873] = 238;
assign img[ 2874] = 238;
assign img[ 2875] = 238;
assign img[ 2876] = 238;
assign img[ 2877] = 238;
assign img[ 2878] = 204;
assign img[ 2879] = 238;
assign img[ 2880] = 238;
assign img[ 2881] = 238;
assign img[ 2882] = 254;
assign img[ 2883] = 255;
assign img[ 2884] = 255;
assign img[ 2885] = 255;
assign img[ 2886] = 238;
assign img[ 2887] = 238;
assign img[ 2888] = 238;
assign img[ 2889] = 207;
assign img[ 2890] = 238;
assign img[ 2891] = 255;
assign img[ 2892] = 255;
assign img[ 2893] = 255;
assign img[ 2894] = 255;
assign img[ 2895] = 255;
assign img[ 2896] = 255;
assign img[ 2897] = 255;
assign img[ 2898] = 223;
assign img[ 2899] = 255;
assign img[ 2900] = 255;
assign img[ 2901] = 239;
assign img[ 2902] = 238;
assign img[ 2903] = 207;
assign img[ 2904] = 255;
assign img[ 2905] = 238;
assign img[ 2906] = 238;
assign img[ 2907] = 206;
assign img[ 2908] = 252;
assign img[ 2909] = 255;
assign img[ 2910] = 255;
assign img[ 2911] = 255;
assign img[ 2912] = 238;
assign img[ 2913] = 238;
assign img[ 2914] = 254;
assign img[ 2915] = 255;
assign img[ 2916] = 255;
assign img[ 2917] = 223;
assign img[ 2918] = 221;
assign img[ 2919] = 253;
assign img[ 2920] = 207;
assign img[ 2921] = 255;
assign img[ 2922] = 239;
assign img[ 2923] = 238;
assign img[ 2924] = 206;
assign img[ 2925] = 238;
assign img[ 2926] = 254;
assign img[ 2927] = 255;
assign img[ 2928] = 221;
assign img[ 2929] = 221;
assign img[ 2930] = 221;
assign img[ 2931] = 221;
assign img[ 2932] = 205;
assign img[ 2933] = 236;
assign img[ 2934] = 254;
assign img[ 2935] = 255;
assign img[ 2936] = 255;
assign img[ 2937] = 255;
assign img[ 2938] = 255;
assign img[ 2939] = 239;
assign img[ 2940] = 238;
assign img[ 2941] = 238;
assign img[ 2942] = 238;
assign img[ 2943] = 238;
assign img[ 2944] = 96;
assign img[ 2945] = 191;
assign img[ 2946] = 251;
assign img[ 2947] = 255;
assign img[ 2948] = 255;
assign img[ 2949] = 255;
assign img[ 2950] = 207;
assign img[ 2951] = 238;
assign img[ 2952] = 238;
assign img[ 2953] = 238;
assign img[ 2954] = 238;
assign img[ 2955] = 255;
assign img[ 2956] = 187;
assign img[ 2957] = 255;
assign img[ 2958] = 255;
assign img[ 2959] = 255;
assign img[ 2960] = 238;
assign img[ 2961] = 254;
assign img[ 2962] = 239;
assign img[ 2963] = 238;
assign img[ 2964] = 238;
assign img[ 2965] = 238;
assign img[ 2966] = 254;
assign img[ 2967] = 255;
assign img[ 2968] = 255;
assign img[ 2969] = 239;
assign img[ 2970] = 170;
assign img[ 2971] = 238;
assign img[ 2972] = 238;
assign img[ 2973] = 255;
assign img[ 2974] = 255;
assign img[ 2975] = 255;
assign img[ 2976] = 155;
assign img[ 2977] = 255;
assign img[ 2978] = 255;
assign img[ 2979] = 255;
assign img[ 2980] = 255;
assign img[ 2981] = 255;
assign img[ 2982] = 255;
assign img[ 2983] = 239;
assign img[ 2984] = 238;
assign img[ 2985] = 255;
assign img[ 2986] = 239;
assign img[ 2987] = 238;
assign img[ 2988] = 238;
assign img[ 2989] = 238;
assign img[ 2990] = 238;
assign img[ 2991] = 238;
assign img[ 2992] = 254;
assign img[ 2993] = 255;
assign img[ 2994] = 255;
assign img[ 2995] = 255;
assign img[ 2996] = 255;
assign img[ 2997] = 255;
assign img[ 2998] = 255;
assign img[ 2999] = 239;
assign img[ 3000] = 238;
assign img[ 3001] = 238;
assign img[ 3002] = 238;
assign img[ 3003] = 238;
assign img[ 3004] = 238;
assign img[ 3005] = 255;
assign img[ 3006] = 238;
assign img[ 3007] = 255;
assign img[ 3008] = 255;
assign img[ 3009] = 255;
assign img[ 3010] = 239;
assign img[ 3011] = 238;
assign img[ 3012] = 238;
assign img[ 3013] = 255;
assign img[ 3014] = 255;
assign img[ 3015] = 255;
assign img[ 3016] = 239;
assign img[ 3017] = 238;
assign img[ 3018] = 238;
assign img[ 3019] = 238;
assign img[ 3020] = 238;
assign img[ 3021] = 238;
assign img[ 3022] = 238;
assign img[ 3023] = 255;
assign img[ 3024] = 255;
assign img[ 3025] = 255;
assign img[ 3026] = 255;
assign img[ 3027] = 255;
assign img[ 3028] = 255;
assign img[ 3029] = 223;
assign img[ 3030] = 255;
assign img[ 3031] = 255;
assign img[ 3032] = 255;
assign img[ 3033] = 255;
assign img[ 3034] = 255;
assign img[ 3035] = 255;
assign img[ 3036] = 255;
assign img[ 3037] = 255;
assign img[ 3038] = 255;
assign img[ 3039] = 223;
assign img[ 3040] = 255;
assign img[ 3041] = 255;
assign img[ 3042] = 255;
assign img[ 3043] = 255;
assign img[ 3044] = 255;
assign img[ 3045] = 255;
assign img[ 3046] = 191;
assign img[ 3047] = 255;
assign img[ 3048] = 255;
assign img[ 3049] = 255;
assign img[ 3050] = 255;
assign img[ 3051] = 239;
assign img[ 3052] = 222;
assign img[ 3053] = 221;
assign img[ 3054] = 236;
assign img[ 3055] = 255;
assign img[ 3056] = 255;
assign img[ 3057] = 255;
assign img[ 3058] = 254;
assign img[ 3059] = 223;
assign img[ 3060] = 221;
assign img[ 3061] = 255;
assign img[ 3062] = 255;
assign img[ 3063] = 255;
assign img[ 3064] = 255;
assign img[ 3065] = 255;
assign img[ 3066] = 238;
assign img[ 3067] = 238;
assign img[ 3068] = 220;
assign img[ 3069] = 255;
assign img[ 3070] = 191;
assign img[ 3071] = 255;
assign img[ 3072] = 96;
assign img[ 3073] = 119;
assign img[ 3074] = 119;
assign img[ 3075] = 255;
assign img[ 3076] = 175;
assign img[ 3077] = 138;
assign img[ 3078] = 136;
assign img[ 3079] = 236;
assign img[ 3080] = 238;
assign img[ 3081] = 239;
assign img[ 3082] = 238;
assign img[ 3083] = 207;
assign img[ 3084] = 204;
assign img[ 3085] = 238;
assign img[ 3086] = 238;
assign img[ 3087] = 255;
assign img[ 3088] = 238;
assign img[ 3089] = 238;
assign img[ 3090] = 238;
assign img[ 3091] = 255;
assign img[ 3092] = 187;
assign img[ 3093] = 255;
assign img[ 3094] = 255;
assign img[ 3095] = 255;
assign img[ 3096] = 255;
assign img[ 3097] = 239;
assign img[ 3098] = 238;
assign img[ 3099] = 238;
assign img[ 3100] = 238;
assign img[ 3101] = 254;
assign img[ 3102] = 255;
assign img[ 3103] = 223;
assign img[ 3104] = 221;
assign img[ 3105] = 255;
assign img[ 3106] = 255;
assign img[ 3107] = 255;
assign img[ 3108] = 255;
assign img[ 3109] = 255;
assign img[ 3110] = 255;
assign img[ 3111] = 223;
assign img[ 3112] = 253;
assign img[ 3113] = 255;
assign img[ 3114] = 175;
assign img[ 3115] = 170;
assign img[ 3116] = 234;
assign img[ 3117] = 238;
assign img[ 3118] = 238;
assign img[ 3119] = 207;
assign img[ 3120] = 238;
assign img[ 3121] = 239;
assign img[ 3122] = 255;
assign img[ 3123] = 255;
assign img[ 3124] = 238;
assign img[ 3125] = 254;
assign img[ 3126] = 238;
assign img[ 3127] = 255;
assign img[ 3128] = 238;
assign img[ 3129] = 255;
assign img[ 3130] = 255;
assign img[ 3131] = 255;
assign img[ 3132] = 255;
assign img[ 3133] = 255;
assign img[ 3134] = 255;
assign img[ 3135] = 255;
assign img[ 3136] = 255;
assign img[ 3137] = 239;
assign img[ 3138] = 238;
assign img[ 3139] = 238;
assign img[ 3140] = 254;
assign img[ 3141] = 239;
assign img[ 3142] = 238;
assign img[ 3143] = 255;
assign img[ 3144] = 255;
assign img[ 3145] = 255;
assign img[ 3146] = 255;
assign img[ 3147] = 255;
assign img[ 3148] = 238;
assign img[ 3149] = 238;
assign img[ 3150] = 238;
assign img[ 3151] = 238;
assign img[ 3152] = 238;
assign img[ 3153] = 238;
assign img[ 3154] = 238;
assign img[ 3155] = 254;
assign img[ 3156] = 255;
assign img[ 3157] = 255;
assign img[ 3158] = 238;
assign img[ 3159] = 238;
assign img[ 3160] = 238;
assign img[ 3161] = 238;
assign img[ 3162] = 238;
assign img[ 3163] = 255;
assign img[ 3164] = 255;
assign img[ 3165] = 255;
assign img[ 3166] = 255;
assign img[ 3167] = 239;
assign img[ 3168] = 206;
assign img[ 3169] = 221;
assign img[ 3170] = 253;
assign img[ 3171] = 255;
assign img[ 3172] = 238;
assign img[ 3173] = 255;
assign img[ 3174] = 223;
assign img[ 3175] = 255;
assign img[ 3176] = 255;
assign img[ 3177] = 239;
assign img[ 3178] = 238;
assign img[ 3179] = 238;
assign img[ 3180] = 238;
assign img[ 3181] = 238;
assign img[ 3182] = 238;
assign img[ 3183] = 238;
assign img[ 3184] = 221;
assign img[ 3185] = 255;
assign img[ 3186] = 254;
assign img[ 3187] = 255;
assign img[ 3188] = 239;
assign img[ 3189] = 255;
assign img[ 3190] = 239;
assign img[ 3191] = 238;
assign img[ 3192] = 238;
assign img[ 3193] = 255;
assign img[ 3194] = 255;
assign img[ 3195] = 255;
assign img[ 3196] = 238;
assign img[ 3197] = 238;
assign img[ 3198] = 238;
assign img[ 3199] = 255;
assign img[ 3200] = 96;
assign img[ 3201] = 238;
assign img[ 3202] = 238;
assign img[ 3203] = 255;
assign img[ 3204] = 255;
assign img[ 3205] = 255;
assign img[ 3206] = 206;
assign img[ 3207] = 238;
assign img[ 3208] = 238;
assign img[ 3209] = 255;
assign img[ 3210] = 255;
assign img[ 3211] = 255;
assign img[ 3212] = 221;
assign img[ 3213] = 221;
assign img[ 3214] = 236;
assign img[ 3215] = 238;
assign img[ 3216] = 220;
assign img[ 3217] = 253;
assign img[ 3218] = 255;
assign img[ 3219] = 255;
assign img[ 3220] = 255;
assign img[ 3221] = 255;
assign img[ 3222] = 255;
assign img[ 3223] = 255;
assign img[ 3224] = 255;
assign img[ 3225] = 255;
assign img[ 3226] = 221;
assign img[ 3227] = 255;
assign img[ 3228] = 255;
assign img[ 3229] = 255;
assign img[ 3230] = 223;
assign img[ 3231] = 221;
assign img[ 3232] = 221;
assign img[ 3233] = 253;
assign img[ 3234] = 255;
assign img[ 3235] = 255;
assign img[ 3236] = 255;
assign img[ 3237] = 239;
assign img[ 3238] = 238;
assign img[ 3239] = 238;
assign img[ 3240] = 238;
assign img[ 3241] = 238;
assign img[ 3242] = 254;
assign img[ 3243] = 223;
assign img[ 3244] = 204;
assign img[ 3245] = 205;
assign img[ 3246] = 236;
assign img[ 3247] = 255;
assign img[ 3248] = 255;
assign img[ 3249] = 255;
assign img[ 3250] = 255;
assign img[ 3251] = 255;
assign img[ 3252] = 255;
assign img[ 3253] = 255;
assign img[ 3254] = 255;
assign img[ 3255] = 255;
assign img[ 3256] = 255;
assign img[ 3257] = 223;
assign img[ 3258] = 204;
assign img[ 3259] = 236;
assign img[ 3260] = 238;
assign img[ 3261] = 206;
assign img[ 3262] = 236;
assign img[ 3263] = 255;
assign img[ 3264] = 255;
assign img[ 3265] = 255;
assign img[ 3266] = 223;
assign img[ 3267] = 255;
assign img[ 3268] = 255;
assign img[ 3269] = 255;
assign img[ 3270] = 205;
assign img[ 3271] = 253;
assign img[ 3272] = 223;
assign img[ 3273] = 253;
assign img[ 3274] = 255;
assign img[ 3275] = 255;
assign img[ 3276] = 255;
assign img[ 3277] = 255;
assign img[ 3278] = 255;
assign img[ 3279] = 255;
assign img[ 3280] = 223;
assign img[ 3281] = 255;
assign img[ 3282] = 239;
assign img[ 3283] = 254;
assign img[ 3284] = 207;
assign img[ 3285] = 204;
assign img[ 3286] = 238;
assign img[ 3287] = 238;
assign img[ 3288] = 254;
assign img[ 3289] = 255;
assign img[ 3290] = 255;
assign img[ 3291] = 255;
assign img[ 3292] = 255;
assign img[ 3293] = 255;
assign img[ 3294] = 255;
assign img[ 3295] = 255;
assign img[ 3296] = 239;
assign img[ 3297] = 255;
assign img[ 3298] = 255;
assign img[ 3299] = 255;
assign img[ 3300] = 255;
assign img[ 3301] = 255;
assign img[ 3302] = 207;
assign img[ 3303] = 238;
assign img[ 3304] = 254;
assign img[ 3305] = 255;
assign img[ 3306] = 255;
assign img[ 3307] = 255;
assign img[ 3308] = 223;
assign img[ 3309] = 255;
assign img[ 3310] = 255;
assign img[ 3311] = 255;
assign img[ 3312] = 255;
assign img[ 3313] = 255;
assign img[ 3314] = 255;
assign img[ 3315] = 207;
assign img[ 3316] = 220;
assign img[ 3317] = 253;
assign img[ 3318] = 255;
assign img[ 3319] = 255;
assign img[ 3320] = 255;
assign img[ 3321] = 223;
assign img[ 3322] = 221;
assign img[ 3323] = 207;
assign img[ 3324] = 204;
assign img[ 3325] = 238;
assign img[ 3326] = 238;
assign img[ 3327] = 238;
assign img[ 3328] = 96;
assign img[ 3329] = 238;
assign img[ 3330] = 238;
assign img[ 3331] = 238;
assign img[ 3332] = 238;
assign img[ 3333] = 238;
assign img[ 3334] = 238;
assign img[ 3335] = 238;
assign img[ 3336] = 238;
assign img[ 3337] = 238;
assign img[ 3338] = 238;
assign img[ 3339] = 222;
assign img[ 3340] = 221;
assign img[ 3341] = 255;
assign img[ 3342] = 223;
assign img[ 3343] = 221;
assign img[ 3344] = 140;
assign img[ 3345] = 186;
assign img[ 3346] = 251;
assign img[ 3347] = 255;
assign img[ 3348] = 255;
assign img[ 3349] = 255;
assign img[ 3350] = 255;
assign img[ 3351] = 255;
assign img[ 3352] = 255;
assign img[ 3353] = 255;
assign img[ 3354] = 239;
assign img[ 3355] = 238;
assign img[ 3356] = 238;
assign img[ 3357] = 238;
assign img[ 3358] = 238;
assign img[ 3359] = 255;
assign img[ 3360] = 239;
assign img[ 3361] = 254;
assign img[ 3362] = 255;
assign img[ 3363] = 255;
assign img[ 3364] = 255;
assign img[ 3365] = 255;
assign img[ 3366] = 238;
assign img[ 3367] = 223;
assign img[ 3368] = 238;
assign img[ 3369] = 238;
assign img[ 3370] = 206;
assign img[ 3371] = 238;
assign img[ 3372] = 238;
assign img[ 3373] = 255;
assign img[ 3374] = 238;
assign img[ 3375] = 238;
assign img[ 3376] = 254;
assign img[ 3377] = 255;
assign img[ 3378] = 255;
assign img[ 3379] = 255;
assign img[ 3380] = 255;
assign img[ 3381] = 255;
assign img[ 3382] = 255;
assign img[ 3383] = 255;
assign img[ 3384] = 255;
assign img[ 3385] = 255;
assign img[ 3386] = 255;
assign img[ 3387] = 255;
assign img[ 3388] = 255;
assign img[ 3389] = 255;
assign img[ 3390] = 255;
assign img[ 3391] = 255;
assign img[ 3392] = 255;
assign img[ 3393] = 255;
assign img[ 3394] = 255;
assign img[ 3395] = 255;
assign img[ 3396] = 255;
assign img[ 3397] = 255;
assign img[ 3398] = 255;
assign img[ 3399] = 239;
assign img[ 3400] = 238;
assign img[ 3401] = 238;
assign img[ 3402] = 254;
assign img[ 3403] = 239;
assign img[ 3404] = 238;
assign img[ 3405] = 238;
assign img[ 3406] = 238;
assign img[ 3407] = 255;
assign img[ 3408] = 255;
assign img[ 3409] = 255;
assign img[ 3410] = 239;
assign img[ 3411] = 238;
assign img[ 3412] = 238;
assign img[ 3413] = 255;
assign img[ 3414] = 255;
assign img[ 3415] = 255;
assign img[ 3416] = 255;
assign img[ 3417] = 255;
assign img[ 3418] = 239;
assign img[ 3419] = 238;
assign img[ 3420] = 254;
assign img[ 3421] = 255;
assign img[ 3422] = 255;
assign img[ 3423] = 255;
assign img[ 3424] = 238;
assign img[ 3425] = 238;
assign img[ 3426] = 238;
assign img[ 3427] = 238;
assign img[ 3428] = 238;
assign img[ 3429] = 255;
assign img[ 3430] = 255;
assign img[ 3431] = 255;
assign img[ 3432] = 255;
assign img[ 3433] = 255;
assign img[ 3434] = 255;
assign img[ 3435] = 255;
assign img[ 3436] = 255;
assign img[ 3437] = 255;
assign img[ 3438] = 255;
assign img[ 3439] = 255;
assign img[ 3440] = 238;
assign img[ 3441] = 222;
assign img[ 3442] = 253;
assign img[ 3443] = 238;
assign img[ 3444] = 238;
assign img[ 3445] = 238;
assign img[ 3446] = 238;
assign img[ 3447] = 238;
assign img[ 3448] = 238;
assign img[ 3449] = 238;
assign img[ 3450] = 238;
assign img[ 3451] = 238;
assign img[ 3452] = 238;
assign img[ 3453] = 238;
assign img[ 3454] = 238;
assign img[ 3455] = 238;
assign img[ 3456] = 80;
assign img[ 3457] = 237;
assign img[ 3458] = 254;
assign img[ 3459] = 239;
assign img[ 3460] = 204;
assign img[ 3461] = 236;
assign img[ 3462] = 174;
assign img[ 3463] = 238;
assign img[ 3464] = 238;
assign img[ 3465] = 238;
assign img[ 3466] = 238;
assign img[ 3467] = 255;
assign img[ 3468] = 221;
assign img[ 3469] = 205;
assign img[ 3470] = 238;
assign img[ 3471] = 238;
assign img[ 3472] = 220;
assign img[ 3473] = 255;
assign img[ 3474] = 255;
assign img[ 3475] = 255;
assign img[ 3476] = 255;
assign img[ 3477] = 255;
assign img[ 3478] = 223;
assign img[ 3479] = 255;
assign img[ 3480] = 255;
assign img[ 3481] = 255;
assign img[ 3482] = 207;
assign img[ 3483] = 238;
assign img[ 3484] = 238;
assign img[ 3485] = 238;
assign img[ 3486] = 238;
assign img[ 3487] = 238;
assign img[ 3488] = 255;
assign img[ 3489] = 255;
assign img[ 3490] = 255;
assign img[ 3491] = 255;
assign img[ 3492] = 255;
assign img[ 3493] = 255;
assign img[ 3494] = 239;
assign img[ 3495] = 239;
assign img[ 3496] = 238;
assign img[ 3497] = 238;
assign img[ 3498] = 238;
assign img[ 3499] = 238;
assign img[ 3500] = 238;
assign img[ 3501] = 238;
assign img[ 3502] = 238;
assign img[ 3503] = 238;
assign img[ 3504] = 254;
assign img[ 3505] = 255;
assign img[ 3506] = 255;
assign img[ 3507] = 254;
assign img[ 3508] = 238;
assign img[ 3509] = 255;
assign img[ 3510] = 255;
assign img[ 3511] = 255;
assign img[ 3512] = 255;
assign img[ 3513] = 255;
assign img[ 3514] = 255;
assign img[ 3515] = 255;
assign img[ 3516] = 255;
assign img[ 3517] = 239;
assign img[ 3518] = 238;
assign img[ 3519] = 255;
assign img[ 3520] = 255;
assign img[ 3521] = 255;
assign img[ 3522] = 255;
assign img[ 3523] = 255;
assign img[ 3524] = 255;
assign img[ 3525] = 255;
assign img[ 3526] = 255;
assign img[ 3527] = 255;
assign img[ 3528] = 221;
assign img[ 3529] = 255;
assign img[ 3530] = 255;
assign img[ 3531] = 255;
assign img[ 3532] = 255;
assign img[ 3533] = 255;
assign img[ 3534] = 255;
assign img[ 3535] = 255;
assign img[ 3536] = 255;
assign img[ 3537] = 255;
assign img[ 3538] = 255;
assign img[ 3539] = 255;
assign img[ 3540] = 255;
assign img[ 3541] = 238;
assign img[ 3542] = 238;
assign img[ 3543] = 238;
assign img[ 3544] = 238;
assign img[ 3545] = 238;
assign img[ 3546] = 238;
assign img[ 3547] = 239;
assign img[ 3548] = 238;
assign img[ 3549] = 255;
assign img[ 3550] = 255;
assign img[ 3551] = 255;
assign img[ 3552] = 255;
assign img[ 3553] = 255;
assign img[ 3554] = 254;
assign img[ 3555] = 255;
assign img[ 3556] = 254;
assign img[ 3557] = 255;
assign img[ 3558] = 221;
assign img[ 3559] = 255;
assign img[ 3560] = 255;
assign img[ 3561] = 255;
assign img[ 3562] = 255;
assign img[ 3563] = 255;
assign img[ 3564] = 207;
assign img[ 3565] = 238;
assign img[ 3566] = 254;
assign img[ 3567] = 255;
assign img[ 3568] = 255;
assign img[ 3569] = 255;
assign img[ 3570] = 239;
assign img[ 3571] = 238;
assign img[ 3572] = 238;
assign img[ 3573] = 254;
assign img[ 3574] = 239;
assign img[ 3575] = 254;
assign img[ 3576] = 254;
assign img[ 3577] = 191;
assign img[ 3578] = 153;
assign img[ 3579] = 171;
assign img[ 3580] = 187;
assign img[ 3581] = 255;
assign img[ 3582] = 255;
assign img[ 3583] = 255;
assign img[ 3584] = 0;
assign img[ 3585] = 128;
assign img[ 3586] = 232;
assign img[ 3587] = 238;
assign img[ 3588] = 238;
assign img[ 3589] = 254;
assign img[ 3590] = 255;
assign img[ 3591] = 255;
assign img[ 3592] = 255;
assign img[ 3593] = 255;
assign img[ 3594] = 255;
assign img[ 3595] = 255;
assign img[ 3596] = 223;
assign img[ 3597] = 221;
assign img[ 3598] = 221;
assign img[ 3599] = 221;
assign img[ 3600] = 204;
assign img[ 3601] = 252;
assign img[ 3602] = 255;
assign img[ 3603] = 255;
assign img[ 3604] = 255;
assign img[ 3605] = 255;
assign img[ 3606] = 239;
assign img[ 3607] = 238;
assign img[ 3608] = 238;
assign img[ 3609] = 207;
assign img[ 3610] = 204;
assign img[ 3611] = 239;
assign img[ 3612] = 238;
assign img[ 3613] = 255;
assign img[ 3614] = 255;
assign img[ 3615] = 255;
assign img[ 3616] = 207;
assign img[ 3617] = 238;
assign img[ 3618] = 238;
assign img[ 3619] = 255;
assign img[ 3620] = 255;
assign img[ 3621] = 255;
assign img[ 3622] = 255;
assign img[ 3623] = 255;
assign img[ 3624] = 255;
assign img[ 3625] = 255;
assign img[ 3626] = 255;
assign img[ 3627] = 255;
assign img[ 3628] = 238;
assign img[ 3629] = 255;
assign img[ 3630] = 255;
assign img[ 3631] = 255;
assign img[ 3632] = 255;
assign img[ 3633] = 255;
assign img[ 3634] = 255;
assign img[ 3635] = 239;
assign img[ 3636] = 238;
assign img[ 3637] = 254;
assign img[ 3638] = 255;
assign img[ 3639] = 254;
assign img[ 3640] = 254;
assign img[ 3641] = 255;
assign img[ 3642] = 255;
assign img[ 3643] = 255;
assign img[ 3644] = 255;
assign img[ 3645] = 255;
assign img[ 3646] = 255;
assign img[ 3647] = 255;
assign img[ 3648] = 255;
assign img[ 3649] = 255;
assign img[ 3650] = 255;
assign img[ 3651] = 255;
assign img[ 3652] = 255;
assign img[ 3653] = 255;
assign img[ 3654] = 255;
assign img[ 3655] = 254;
assign img[ 3656] = 255;
assign img[ 3657] = 255;
assign img[ 3658] = 255;
assign img[ 3659] = 223;
assign img[ 3660] = 221;
assign img[ 3661] = 255;
assign img[ 3662] = 255;
assign img[ 3663] = 255;
assign img[ 3664] = 239;
assign img[ 3665] = 238;
assign img[ 3666] = 206;
assign img[ 3667] = 238;
assign img[ 3668] = 238;
assign img[ 3669] = 254;
assign img[ 3670] = 255;
assign img[ 3671] = 255;
assign img[ 3672] = 255;
assign img[ 3673] = 255;
assign img[ 3674] = 255;
assign img[ 3675] = 239;
assign img[ 3676] = 254;
assign img[ 3677] = 255;
assign img[ 3678] = 255;
assign img[ 3679] = 223;
assign img[ 3680] = 236;
assign img[ 3681] = 223;
assign img[ 3682] = 253;
assign img[ 3683] = 255;
assign img[ 3684] = 255;
assign img[ 3685] = 255;
assign img[ 3686] = 239;
assign img[ 3687] = 255;
assign img[ 3688] = 255;
assign img[ 3689] = 255;
assign img[ 3690] = 255;
assign img[ 3691] = 255;
assign img[ 3692] = 255;
assign img[ 3693] = 255;
assign img[ 3694] = 255;
assign img[ 3695] = 255;
assign img[ 3696] = 204;
assign img[ 3697] = 204;
assign img[ 3698] = 204;
assign img[ 3699] = 206;
assign img[ 3700] = 204;
assign img[ 3701] = 238;
assign img[ 3702] = 238;
assign img[ 3703] = 238;
assign img[ 3704] = 238;
assign img[ 3705] = 255;
assign img[ 3706] = 255;
assign img[ 3707] = 223;
assign img[ 3708] = 221;
assign img[ 3709] = 253;
assign img[ 3710] = 223;
assign img[ 3711] = 221;
assign img[ 3712] = 96;
assign img[ 3713] = 223;
assign img[ 3714] = 221;
assign img[ 3715] = 153;
assign img[ 3716] = 249;
assign img[ 3717] = 255;
assign img[ 3718] = 207;
assign img[ 3719] = 238;
assign img[ 3720] = 238;
assign img[ 3721] = 238;
assign img[ 3722] = 254;
assign img[ 3723] = 207;
assign img[ 3724] = 204;
assign img[ 3725] = 238;
assign img[ 3726] = 238;
assign img[ 3727] = 238;
assign img[ 3728] = 204;
assign img[ 3729] = 204;
assign img[ 3730] = 236;
assign img[ 3731] = 206;
assign img[ 3732] = 236;
assign img[ 3733] = 238;
assign img[ 3734] = 238;
assign img[ 3735] = 255;
assign img[ 3736] = 255;
assign img[ 3737] = 255;
assign img[ 3738] = 255;
assign img[ 3739] = 238;
assign img[ 3740] = 255;
assign img[ 3741] = 255;
assign img[ 3742] = 223;
assign img[ 3743] = 157;
assign img[ 3744] = 153;
assign img[ 3745] = 253;
assign img[ 3746] = 255;
assign img[ 3747] = 255;
assign img[ 3748] = 255;
assign img[ 3749] = 255;
assign img[ 3750] = 255;
assign img[ 3751] = 255;
assign img[ 3752] = 255;
assign img[ 3753] = 255;
assign img[ 3754] = 239;
assign img[ 3755] = 238;
assign img[ 3756] = 255;
assign img[ 3757] = 255;
assign img[ 3758] = 255;
assign img[ 3759] = 255;
assign img[ 3760] = 255;
assign img[ 3761] = 255;
assign img[ 3762] = 255;
assign img[ 3763] = 255;
assign img[ 3764] = 238;
assign img[ 3765] = 238;
assign img[ 3766] = 190;
assign img[ 3767] = 255;
assign img[ 3768] = 255;
assign img[ 3769] = 255;
assign img[ 3770] = 223;
assign img[ 3771] = 255;
assign img[ 3772] = 255;
assign img[ 3773] = 255;
assign img[ 3774] = 255;
assign img[ 3775] = 255;
assign img[ 3776] = 255;
assign img[ 3777] = 255;
assign img[ 3778] = 255;
assign img[ 3779] = 255;
assign img[ 3780] = 255;
assign img[ 3781] = 255;
assign img[ 3782] = 255;
assign img[ 3783] = 255;
assign img[ 3784] = 255;
assign img[ 3785] = 255;
assign img[ 3786] = 255;
assign img[ 3787] = 239;
assign img[ 3788] = 238;
assign img[ 3789] = 238;
assign img[ 3790] = 254;
assign img[ 3791] = 255;
assign img[ 3792] = 255;
assign img[ 3793] = 255;
assign img[ 3794] = 255;
assign img[ 3795] = 255;
assign img[ 3796] = 255;
assign img[ 3797] = 255;
assign img[ 3798] = 255;
assign img[ 3799] = 255;
assign img[ 3800] = 255;
assign img[ 3801] = 255;
assign img[ 3802] = 255;
assign img[ 3803] = 255;
assign img[ 3804] = 255;
assign img[ 3805] = 255;
assign img[ 3806] = 255;
assign img[ 3807] = 223;
assign img[ 3808] = 221;
assign img[ 3809] = 221;
assign img[ 3810] = 255;
assign img[ 3811] = 255;
assign img[ 3812] = 255;
assign img[ 3813] = 239;
assign img[ 3814] = 254;
assign img[ 3815] = 255;
assign img[ 3816] = 255;
assign img[ 3817] = 239;
assign img[ 3818] = 238;
assign img[ 3819] = 255;
assign img[ 3820] = 255;
assign img[ 3821] = 255;
assign img[ 3822] = 255;
assign img[ 3823] = 223;
assign img[ 3824] = 221;
assign img[ 3825] = 253;
assign img[ 3826] = 255;
assign img[ 3827] = 239;
assign img[ 3828] = 206;
assign img[ 3829] = 221;
assign img[ 3830] = 253;
assign img[ 3831] = 255;
assign img[ 3832] = 255;
assign img[ 3833] = 223;
assign img[ 3834] = 221;
assign img[ 3835] = 221;
assign img[ 3836] = 157;
assign img[ 3837] = 153;
assign img[ 3838] = 153;
assign img[ 3839] = 255;
assign img[ 3840] = 112;
assign img[ 3841] = 255;
assign img[ 3842] = 255;
assign img[ 3843] = 223;
assign img[ 3844] = 221;
assign img[ 3845] = 255;
assign img[ 3846] = 174;
assign img[ 3847] = 238;
assign img[ 3848] = 238;
assign img[ 3849] = 255;
assign img[ 3850] = 238;
assign img[ 3851] = 255;
assign img[ 3852] = 221;
assign img[ 3853] = 255;
assign img[ 3854] = 255;
assign img[ 3855] = 255;
assign img[ 3856] = 238;
assign img[ 3857] = 238;
assign img[ 3858] = 255;
assign img[ 3859] = 255;
assign img[ 3860] = 255;
assign img[ 3861] = 255;
assign img[ 3862] = 255;
assign img[ 3863] = 255;
assign img[ 3864] = 255;
assign img[ 3865] = 207;
assign img[ 3866] = 204;
assign img[ 3867] = 238;
assign img[ 3868] = 238;
assign img[ 3869] = 255;
assign img[ 3870] = 255;
assign img[ 3871] = 175;
assign img[ 3872] = 202;
assign img[ 3873] = 255;
assign img[ 3874] = 223;
assign img[ 3875] = 255;
assign img[ 3876] = 255;
assign img[ 3877] = 255;
assign img[ 3878] = 238;
assign img[ 3879] = 255;
assign img[ 3880] = 238;
assign img[ 3881] = 238;
assign img[ 3882] = 238;
assign img[ 3883] = 238;
assign img[ 3884] = 170;
assign img[ 3885] = 254;
assign img[ 3886] = 254;
assign img[ 3887] = 255;
assign img[ 3888] = 255;
assign img[ 3889] = 255;
assign img[ 3890] = 255;
assign img[ 3891] = 255;
assign img[ 3892] = 255;
assign img[ 3893] = 255;
assign img[ 3894] = 255;
assign img[ 3895] = 255;
assign img[ 3896] = 255;
assign img[ 3897] = 255;
assign img[ 3898] = 255;
assign img[ 3899] = 255;
assign img[ 3900] = 255;
assign img[ 3901] = 255;
assign img[ 3902] = 221;
assign img[ 3903] = 255;
assign img[ 3904] = 255;
assign img[ 3905] = 255;
assign img[ 3906] = 255;
assign img[ 3907] = 255;
assign img[ 3908] = 255;
assign img[ 3909] = 239;
assign img[ 3910] = 238;
assign img[ 3911] = 238;
assign img[ 3912] = 254;
assign img[ 3913] = 255;
assign img[ 3914] = 255;
assign img[ 3915] = 255;
assign img[ 3916] = 206;
assign img[ 3917] = 238;
assign img[ 3918] = 238;
assign img[ 3919] = 255;
assign img[ 3920] = 255;
assign img[ 3921] = 255;
assign img[ 3922] = 255;
assign img[ 3923] = 255;
assign img[ 3924] = 255;
assign img[ 3925] = 255;
assign img[ 3926] = 255;
assign img[ 3927] = 255;
assign img[ 3928] = 255;
assign img[ 3929] = 255;
assign img[ 3930] = 239;
assign img[ 3931] = 238;
assign img[ 3932] = 238;
assign img[ 3933] = 238;
assign img[ 3934] = 254;
assign img[ 3935] = 223;
assign img[ 3936] = 157;
assign img[ 3937] = 187;
assign img[ 3938] = 251;
assign img[ 3939] = 255;
assign img[ 3940] = 255;
assign img[ 3941] = 255;
assign img[ 3942] = 223;
assign img[ 3943] = 255;
assign img[ 3944] = 255;
assign img[ 3945] = 255;
assign img[ 3946] = 255;
assign img[ 3947] = 255;
assign img[ 3948] = 223;
assign img[ 3949] = 255;
assign img[ 3950] = 255;
assign img[ 3951] = 255;
assign img[ 3952] = 239;
assign img[ 3953] = 238;
assign img[ 3954] = 238;
assign img[ 3955] = 255;
assign img[ 3956] = 239;
assign img[ 3957] = 238;
assign img[ 3958] = 238;
assign img[ 3959] = 238;
assign img[ 3960] = 238;
assign img[ 3961] = 255;
assign img[ 3962] = 239;
assign img[ 3963] = 238;
assign img[ 3964] = 238;
assign img[ 3965] = 255;
assign img[ 3966] = 255;
assign img[ 3967] = 255;
assign img[ 3968] = 96;
assign img[ 3969] = 238;
assign img[ 3970] = 238;
assign img[ 3971] = 206;
assign img[ 3972] = 204;
assign img[ 3973] = 236;
assign img[ 3974] = 254;
assign img[ 3975] = 255;
assign img[ 3976] = 255;
assign img[ 3977] = 255;
assign img[ 3978] = 238;
assign img[ 3979] = 238;
assign img[ 3980] = 238;
assign img[ 3981] = 238;
assign img[ 3982] = 238;
assign img[ 3983] = 238;
assign img[ 3984] = 204;
assign img[ 3985] = 204;
assign img[ 3986] = 236;
assign img[ 3987] = 223;
assign img[ 3988] = 204;
assign img[ 3989] = 238;
assign img[ 3990] = 238;
assign img[ 3991] = 238;
assign img[ 3992] = 238;
assign img[ 3993] = 191;
assign img[ 3994] = 171;
assign img[ 3995] = 238;
assign img[ 3996] = 238;
assign img[ 3997] = 238;
assign img[ 3998] = 254;
assign img[ 3999] = 239;
assign img[ 4000] = 238;
assign img[ 4001] = 238;
assign img[ 4002] = 238;
assign img[ 4003] = 255;
assign img[ 4004] = 191;
assign img[ 4005] = 255;
assign img[ 4006] = 255;
assign img[ 4007] = 255;
assign img[ 4008] = 255;
assign img[ 4009] = 255;
assign img[ 4010] = 239;
assign img[ 4011] = 238;
assign img[ 4012] = 254;
assign img[ 4013] = 223;
assign img[ 4014] = 255;
assign img[ 4015] = 255;
assign img[ 4016] = 255;
assign img[ 4017] = 255;
assign img[ 4018] = 255;
assign img[ 4019] = 255;
assign img[ 4020] = 255;
assign img[ 4021] = 255;
assign img[ 4022] = 239;
assign img[ 4023] = 238;
assign img[ 4024] = 238;
assign img[ 4025] = 255;
assign img[ 4026] = 223;
assign img[ 4027] = 255;
assign img[ 4028] = 255;
assign img[ 4029] = 255;
assign img[ 4030] = 255;
assign img[ 4031] = 255;
assign img[ 4032] = 255;
assign img[ 4033] = 255;
assign img[ 4034] = 255;
assign img[ 4035] = 255;
assign img[ 4036] = 255;
assign img[ 4037] = 223;
assign img[ 4038] = 255;
assign img[ 4039] = 255;
assign img[ 4040] = 255;
assign img[ 4041] = 255;
assign img[ 4042] = 255;
assign img[ 4043] = 255;
assign img[ 4044] = 255;
assign img[ 4045] = 255;
assign img[ 4046] = 255;
assign img[ 4047] = 255;
assign img[ 4048] = 239;
assign img[ 4049] = 238;
assign img[ 4050] = 222;
assign img[ 4051] = 205;
assign img[ 4052] = 220;
assign img[ 4053] = 221;
assign img[ 4054] = 236;
assign img[ 4055] = 238;
assign img[ 4056] = 238;
assign img[ 4057] = 254;
assign img[ 4058] = 238;
assign img[ 4059] = 255;
assign img[ 4060] = 255;
assign img[ 4061] = 255;
assign img[ 4062] = 255;
assign img[ 4063] = 239;
assign img[ 4064] = 238;
assign img[ 4065] = 254;
assign img[ 4066] = 255;
assign img[ 4067] = 255;
assign img[ 4068] = 254;
assign img[ 4069] = 255;
assign img[ 4070] = 238;
assign img[ 4071] = 238;
assign img[ 4072] = 254;
assign img[ 4073] = 255;
assign img[ 4074] = 238;
assign img[ 4075] = 255;
assign img[ 4076] = 238;
assign img[ 4077] = 238;
assign img[ 4078] = 254;
assign img[ 4079] = 239;
assign img[ 4080] = 220;
assign img[ 4081] = 253;
assign img[ 4082] = 255;
assign img[ 4083] = 255;
assign img[ 4084] = 255;
assign img[ 4085] = 255;
assign img[ 4086] = 255;
assign img[ 4087] = 255;
assign img[ 4088] = 255;
assign img[ 4089] = 223;
assign img[ 4090] = 221;
assign img[ 4091] = 223;
assign img[ 4092] = 221;
assign img[ 4093] = 253;
assign img[ 4094] = 255;
assign img[ 4095] = 255;
assign img[ 4096] = 96;
assign img[ 4097] = 206;
assign img[ 4098] = 252;
assign img[ 4099] = 255;
assign img[ 4100] = 205;
assign img[ 4101] = 238;
assign img[ 4102] = 238;
assign img[ 4103] = 238;
assign img[ 4104] = 238;
assign img[ 4105] = 238;
assign img[ 4106] = 238;
assign img[ 4107] = 222;
assign img[ 4108] = 253;
assign img[ 4109] = 255;
assign img[ 4110] = 255;
assign img[ 4111] = 238;
assign img[ 4112] = 238;
assign img[ 4113] = 238;
assign img[ 4114] = 254;
assign img[ 4115] = 223;
assign img[ 4116] = 238;
assign img[ 4117] = 238;
assign img[ 4118] = 254;
assign img[ 4119] = 255;
assign img[ 4120] = 255;
assign img[ 4121] = 191;
assign img[ 4122] = 170;
assign img[ 4123] = 238;
assign img[ 4124] = 254;
assign img[ 4125] = 255;
assign img[ 4126] = 255;
assign img[ 4127] = 207;
assign img[ 4128] = 136;
assign img[ 4129] = 238;
assign img[ 4130] = 238;
assign img[ 4131] = 255;
assign img[ 4132] = 255;
assign img[ 4133] = 255;
assign img[ 4134] = 255;
assign img[ 4135] = 255;
assign img[ 4136] = 255;
assign img[ 4137] = 255;
assign img[ 4138] = 239;
assign img[ 4139] = 238;
assign img[ 4140] = 238;
assign img[ 4141] = 238;
assign img[ 4142] = 238;
assign img[ 4143] = 238;
assign img[ 4144] = 255;
assign img[ 4145] = 255;
assign img[ 4146] = 255;
assign img[ 4147] = 255;
assign img[ 4148] = 238;
assign img[ 4149] = 238;
assign img[ 4150] = 238;
assign img[ 4151] = 254;
assign img[ 4152] = 254;
assign img[ 4153] = 255;
assign img[ 4154] = 255;
assign img[ 4155] = 255;
assign img[ 4156] = 255;
assign img[ 4157] = 223;
assign img[ 4158] = 255;
assign img[ 4159] = 255;
assign img[ 4160] = 255;
assign img[ 4161] = 255;
assign img[ 4162] = 255;
assign img[ 4163] = 255;
assign img[ 4164] = 255;
assign img[ 4165] = 239;
assign img[ 4166] = 238;
assign img[ 4167] = 223;
assign img[ 4168] = 253;
assign img[ 4169] = 255;
assign img[ 4170] = 255;
assign img[ 4171] = 223;
assign img[ 4172] = 239;
assign img[ 4173] = 238;
assign img[ 4174] = 238;
assign img[ 4175] = 255;
assign img[ 4176] = 255;
assign img[ 4177] = 255;
assign img[ 4178] = 255;
assign img[ 4179] = 223;
assign img[ 4180] = 253;
assign img[ 4181] = 255;
assign img[ 4182] = 238;
assign img[ 4183] = 255;
assign img[ 4184] = 255;
assign img[ 4185] = 255;
assign img[ 4186] = 223;
assign img[ 4187] = 221;
assign img[ 4188] = 253;
assign img[ 4189] = 255;
assign img[ 4190] = 255;
assign img[ 4191] = 255;
assign img[ 4192] = 223;
assign img[ 4193] = 221;
assign img[ 4194] = 253;
assign img[ 4195] = 255;
assign img[ 4196] = 255;
assign img[ 4197] = 255;
assign img[ 4198] = 238;
assign img[ 4199] = 238;
assign img[ 4200] = 238;
assign img[ 4201] = 238;
assign img[ 4202] = 238;
assign img[ 4203] = 238;
assign img[ 4204] = 206;
assign img[ 4205] = 254;
assign img[ 4206] = 255;
assign img[ 4207] = 255;
assign img[ 4208] = 255;
assign img[ 4209] = 255;
assign img[ 4210] = 255;
assign img[ 4211] = 255;
assign img[ 4212] = 238;
assign img[ 4213] = 239;
assign img[ 4214] = 238;
assign img[ 4215] = 238;
assign img[ 4216] = 238;
assign img[ 4217] = 238;
assign img[ 4218] = 238;
assign img[ 4219] = 255;
assign img[ 4220] = 205;
assign img[ 4221] = 254;
assign img[ 4222] = 223;
assign img[ 4223] = 255;
assign img[ 4224] = 96;
assign img[ 4225] = 239;
assign img[ 4226] = 238;
assign img[ 4227] = 238;
assign img[ 4228] = 206;
assign img[ 4229] = 238;
assign img[ 4230] = 255;
assign img[ 4231] = 255;
assign img[ 4232] = 255;
assign img[ 4233] = 255;
assign img[ 4234] = 239;
assign img[ 4235] = 238;
assign img[ 4236] = 238;
assign img[ 4237] = 254;
assign img[ 4238] = 191;
assign img[ 4239] = 171;
assign img[ 4240] = 200;
assign img[ 4241] = 252;
assign img[ 4242] = 255;
assign img[ 4243] = 255;
assign img[ 4244] = 255;
assign img[ 4245] = 255;
assign img[ 4246] = 223;
assign img[ 4247] = 255;
assign img[ 4248] = 255;
assign img[ 4249] = 255;
assign img[ 4250] = 238;
assign img[ 4251] = 238;
assign img[ 4252] = 238;
assign img[ 4253] = 255;
assign img[ 4254] = 255;
assign img[ 4255] = 223;
assign img[ 4256] = 221;
assign img[ 4257] = 253;
assign img[ 4258] = 254;
assign img[ 4259] = 255;
assign img[ 4260] = 255;
assign img[ 4261] = 255;
assign img[ 4262] = 255;
assign img[ 4263] = 255;
assign img[ 4264] = 255;
assign img[ 4265] = 255;
assign img[ 4266] = 239;
assign img[ 4267] = 238;
assign img[ 4268] = 238;
assign img[ 4269] = 238;
assign img[ 4270] = 238;
assign img[ 4271] = 238;
assign img[ 4272] = 254;
assign img[ 4273] = 255;
assign img[ 4274] = 255;
assign img[ 4275] = 239;
assign img[ 4276] = 238;
assign img[ 4277] = 255;
assign img[ 4278] = 255;
assign img[ 4279] = 255;
assign img[ 4280] = 255;
assign img[ 4281] = 255;
assign img[ 4282] = 255;
assign img[ 4283] = 223;
assign img[ 4284] = 253;
assign img[ 4285] = 223;
assign img[ 4286] = 253;
assign img[ 4287] = 255;
assign img[ 4288] = 255;
assign img[ 4289] = 255;
assign img[ 4290] = 255;
assign img[ 4291] = 255;
assign img[ 4292] = 255;
assign img[ 4293] = 255;
assign img[ 4294] = 255;
assign img[ 4295] = 255;
assign img[ 4296] = 255;
assign img[ 4297] = 255;
assign img[ 4298] = 255;
assign img[ 4299] = 255;
assign img[ 4300] = 255;
assign img[ 4301] = 255;
assign img[ 4302] = 255;
assign img[ 4303] = 255;
assign img[ 4304] = 255;
assign img[ 4305] = 255;
assign img[ 4306] = 255;
assign img[ 4307] = 255;
assign img[ 4308] = 255;
assign img[ 4309] = 255;
assign img[ 4310] = 206;
assign img[ 4311] = 238;
assign img[ 4312] = 254;
assign img[ 4313] = 255;
assign img[ 4314] = 239;
assign img[ 4315] = 255;
assign img[ 4316] = 255;
assign img[ 4317] = 255;
assign img[ 4318] = 255;
assign img[ 4319] = 191;
assign img[ 4320] = 255;
assign img[ 4321] = 255;
assign img[ 4322] = 255;
assign img[ 4323] = 255;
assign img[ 4324] = 255;
assign img[ 4325] = 255;
assign img[ 4326] = 204;
assign img[ 4327] = 236;
assign img[ 4328] = 254;
assign img[ 4329] = 223;
assign img[ 4330] = 221;
assign img[ 4331] = 255;
assign img[ 4332] = 255;
assign img[ 4333] = 255;
assign img[ 4334] = 255;
assign img[ 4335] = 255;
assign img[ 4336] = 221;
assign img[ 4337] = 173;
assign img[ 4338] = 136;
assign img[ 4339] = 255;
assign img[ 4340] = 221;
assign img[ 4341] = 239;
assign img[ 4342] = 238;
assign img[ 4343] = 238;
assign img[ 4344] = 238;
assign img[ 4345] = 255;
assign img[ 4346] = 255;
assign img[ 4347] = 239;
assign img[ 4348] = 220;
assign img[ 4349] = 255;
assign img[ 4350] = 239;
assign img[ 4351] = 238;
assign img[ 4352] = 96;
assign img[ 4353] = 239;
assign img[ 4354] = 255;
assign img[ 4355] = 207;
assign img[ 4356] = 172;
assign img[ 4357] = 138;
assign img[ 4358] = 200;
assign img[ 4359] = 236;
assign img[ 4360] = 238;
assign img[ 4361] = 254;
assign img[ 4362] = 238;
assign img[ 4363] = 238;
assign img[ 4364] = 238;
assign img[ 4365] = 255;
assign img[ 4366] = 255;
assign img[ 4367] = 223;
assign img[ 4368] = 221;
assign img[ 4369] = 255;
assign img[ 4370] = 255;
assign img[ 4371] = 223;
assign img[ 4372] = 236;
assign img[ 4373] = 238;
assign img[ 4374] = 255;
assign img[ 4375] = 255;
assign img[ 4376] = 255;
assign img[ 4377] = 239;
assign img[ 4378] = 238;
assign img[ 4379] = 238;
assign img[ 4380] = 238;
assign img[ 4381] = 254;
assign img[ 4382] = 239;
assign img[ 4383] = 239;
assign img[ 4384] = 204;
assign img[ 4385] = 236;
assign img[ 4386] = 238;
assign img[ 4387] = 255;
assign img[ 4388] = 255;
assign img[ 4389] = 255;
assign img[ 4390] = 255;
assign img[ 4391] = 255;
assign img[ 4392] = 255;
assign img[ 4393] = 255;
assign img[ 4394] = 255;
assign img[ 4395] = 255;
assign img[ 4396] = 206;
assign img[ 4397] = 204;
assign img[ 4398] = 236;
assign img[ 4399] = 223;
assign img[ 4400] = 253;
assign img[ 4401] = 255;
assign img[ 4402] = 255;
assign img[ 4403] = 255;
assign img[ 4404] = 239;
assign img[ 4405] = 238;
assign img[ 4406] = 238;
assign img[ 4407] = 238;
assign img[ 4408] = 238;
assign img[ 4409] = 254;
assign img[ 4410] = 238;
assign img[ 4411] = 255;
assign img[ 4412] = 254;
assign img[ 4413] = 191;
assign img[ 4414] = 255;
assign img[ 4415] = 255;
assign img[ 4416] = 255;
assign img[ 4417] = 255;
assign img[ 4418] = 255;
assign img[ 4419] = 255;
assign img[ 4420] = 223;
assign img[ 4421] = 223;
assign img[ 4422] = 255;
assign img[ 4423] = 239;
assign img[ 4424] = 238;
assign img[ 4425] = 238;
assign img[ 4426] = 238;
assign img[ 4427] = 255;
assign img[ 4428] = 238;
assign img[ 4429] = 238;
assign img[ 4430] = 238;
assign img[ 4431] = 255;
assign img[ 4432] = 255;
assign img[ 4433] = 255;
assign img[ 4434] = 255;
assign img[ 4435] = 223;
assign img[ 4436] = 236;
assign img[ 4437] = 238;
assign img[ 4438] = 254;
assign img[ 4439] = 255;
assign img[ 4440] = 191;
assign img[ 4441] = 255;
assign img[ 4442] = 255;
assign img[ 4443] = 255;
assign img[ 4444] = 255;
assign img[ 4445] = 255;
assign img[ 4446] = 255;
assign img[ 4447] = 239;
assign img[ 4448] = 238;
assign img[ 4449] = 223;
assign img[ 4450] = 253;
assign img[ 4451] = 255;
assign img[ 4452] = 238;
assign img[ 4453] = 223;
assign img[ 4454] = 221;
assign img[ 4455] = 253;
assign img[ 4456] = 238;
assign img[ 4457] = 239;
assign img[ 4458] = 238;
assign img[ 4459] = 238;
assign img[ 4460] = 206;
assign img[ 4461] = 238;
assign img[ 4462] = 238;
assign img[ 4463] = 255;
assign img[ 4464] = 255;
assign img[ 4465] = 255;
assign img[ 4466] = 255;
assign img[ 4467] = 255;
assign img[ 4468] = 207;
assign img[ 4469] = 205;
assign img[ 4470] = 221;
assign img[ 4471] = 255;
assign img[ 4472] = 255;
assign img[ 4473] = 239;
assign img[ 4474] = 254;
assign img[ 4475] = 239;
assign img[ 4476] = 206;
assign img[ 4477] = 255;
assign img[ 4478] = 239;
assign img[ 4479] = 238;
assign img[ 4480] = 96;
assign img[ 4481] = 238;
assign img[ 4482] = 238;
assign img[ 4483] = 223;
assign img[ 4484] = 221;
assign img[ 4485] = 253;
assign img[ 4486] = 204;
assign img[ 4487] = 236;
assign img[ 4488] = 238;
assign img[ 4489] = 238;
assign img[ 4490] = 238;
assign img[ 4491] = 223;
assign img[ 4492] = 236;
assign img[ 4493] = 238;
assign img[ 4494] = 254;
assign img[ 4495] = 255;
assign img[ 4496] = 255;
assign img[ 4497] = 255;
assign img[ 4498] = 255;
assign img[ 4499] = 223;
assign img[ 4500] = 253;
assign img[ 4501] = 238;
assign img[ 4502] = 238;
assign img[ 4503] = 254;
assign img[ 4504] = 255;
assign img[ 4505] = 255;
assign img[ 4506] = 255;
assign img[ 4507] = 255;
assign img[ 4508] = 255;
assign img[ 4509] = 255;
assign img[ 4510] = 255;
assign img[ 4511] = 223;
assign img[ 4512] = 204;
assign img[ 4513] = 236;
assign img[ 4514] = 238;
assign img[ 4515] = 238;
assign img[ 4516] = 238;
assign img[ 4517] = 238;
assign img[ 4518] = 238;
assign img[ 4519] = 255;
assign img[ 4520] = 255;
assign img[ 4521] = 255;
assign img[ 4522] = 255;
assign img[ 4523] = 255;
assign img[ 4524] = 255;
assign img[ 4525] = 223;
assign img[ 4526] = 253;
assign img[ 4527] = 255;
assign img[ 4528] = 255;
assign img[ 4529] = 255;
assign img[ 4530] = 255;
assign img[ 4531] = 255;
assign img[ 4532] = 255;
assign img[ 4533] = 255;
assign img[ 4534] = 255;
assign img[ 4535] = 255;
assign img[ 4536] = 255;
assign img[ 4537] = 255;
assign img[ 4538] = 255;
assign img[ 4539] = 255;
assign img[ 4540] = 255;
assign img[ 4541] = 255;
assign img[ 4542] = 221;
assign img[ 4543] = 255;
assign img[ 4544] = 255;
assign img[ 4545] = 255;
assign img[ 4546] = 255;
assign img[ 4547] = 255;
assign img[ 4548] = 255;
assign img[ 4549] = 255;
assign img[ 4550] = 255;
assign img[ 4551] = 255;
assign img[ 4552] = 255;
assign img[ 4553] = 255;
assign img[ 4554] = 255;
assign img[ 4555] = 255;
assign img[ 4556] = 255;
assign img[ 4557] = 239;
assign img[ 4558] = 238;
assign img[ 4559] = 255;
assign img[ 4560] = 239;
assign img[ 4561] = 238;
assign img[ 4562] = 222;
assign img[ 4563] = 221;
assign img[ 4564] = 253;
assign img[ 4565] = 255;
assign img[ 4566] = 255;
assign img[ 4567] = 255;
assign img[ 4568] = 255;
assign img[ 4569] = 255;
assign img[ 4570] = 255;
assign img[ 4571] = 239;
assign img[ 4572] = 238;
assign img[ 4573] = 238;
assign img[ 4574] = 238;
assign img[ 4575] = 206;
assign img[ 4576] = 204;
assign img[ 4577] = 236;
assign img[ 4578] = 254;
assign img[ 4579] = 255;
assign img[ 4580] = 238;
assign img[ 4581] = 238;
assign img[ 4582] = 238;
assign img[ 4583] = 238;
assign img[ 4584] = 254;
assign img[ 4585] = 255;
assign img[ 4586] = 238;
assign img[ 4587] = 238;
assign img[ 4588] = 206;
assign img[ 4589] = 204;
assign img[ 4590] = 252;
assign img[ 4591] = 239;
assign img[ 4592] = 220;
assign img[ 4593] = 253;
assign img[ 4594] = 255;
assign img[ 4595] = 255;
assign img[ 4596] = 255;
assign img[ 4597] = 255;
assign img[ 4598] = 255;
assign img[ 4599] = 255;
assign img[ 4600] = 255;
assign img[ 4601] = 255;
assign img[ 4602] = 221;
assign img[ 4603] = 221;
assign img[ 4604] = 221;
assign img[ 4605] = 253;
assign img[ 4606] = 255;
assign img[ 4607] = 255;
assign img[ 4608] = 96;
assign img[ 4609] = 238;
assign img[ 4610] = 254;
assign img[ 4611] = 255;
assign img[ 4612] = 223;
assign img[ 4613] = 221;
assign img[ 4614] = 204;
assign img[ 4615] = 220;
assign img[ 4616] = 253;
assign img[ 4617] = 255;
assign img[ 4618] = 255;
assign img[ 4619] = 239;
assign img[ 4620] = 238;
assign img[ 4621] = 238;
assign img[ 4622] = 238;
assign img[ 4623] = 238;
assign img[ 4624] = 238;
assign img[ 4625] = 238;
assign img[ 4626] = 254;
assign img[ 4627] = 255;
assign img[ 4628] = 255;
assign img[ 4629] = 255;
assign img[ 4630] = 239;
assign img[ 4631] = 238;
assign img[ 4632] = 238;
assign img[ 4633] = 207;
assign img[ 4634] = 204;
assign img[ 4635] = 238;
assign img[ 4636] = 238;
assign img[ 4637] = 255;
assign img[ 4638] = 255;
assign img[ 4639] = 191;
assign img[ 4640] = 251;
assign img[ 4641] = 255;
assign img[ 4642] = 191;
assign img[ 4643] = 255;
assign img[ 4644] = 255;
assign img[ 4645] = 255;
assign img[ 4646] = 255;
assign img[ 4647] = 239;
assign img[ 4648] = 238;
assign img[ 4649] = 238;
assign img[ 4650] = 222;
assign img[ 4651] = 255;
assign img[ 4652] = 255;
assign img[ 4653] = 255;
assign img[ 4654] = 255;
assign img[ 4655] = 255;
assign img[ 4656] = 255;
assign img[ 4657] = 255;
assign img[ 4658] = 255;
assign img[ 4659] = 255;
assign img[ 4660] = 255;
assign img[ 4661] = 255;
assign img[ 4662] = 255;
assign img[ 4663] = 255;
assign img[ 4664] = 255;
assign img[ 4665] = 255;
assign img[ 4666] = 222;
assign img[ 4667] = 255;
assign img[ 4668] = 223;
assign img[ 4669] = 157;
assign img[ 4670] = 248;
assign img[ 4671] = 255;
assign img[ 4672] = 255;
assign img[ 4673] = 255;
assign img[ 4674] = 191;
assign img[ 4675] = 139;
assign img[ 4676] = 232;
assign img[ 4677] = 255;
assign img[ 4678] = 255;
assign img[ 4679] = 255;
assign img[ 4680] = 255;
assign img[ 4681] = 255;
assign img[ 4682] = 255;
assign img[ 4683] = 255;
assign img[ 4684] = 255;
assign img[ 4685] = 255;
assign img[ 4686] = 238;
assign img[ 4687] = 255;
assign img[ 4688] = 255;
assign img[ 4689] = 255;
assign img[ 4690] = 223;
assign img[ 4691] = 255;
assign img[ 4692] = 255;
assign img[ 4693] = 255;
assign img[ 4694] = 255;
assign img[ 4695] = 255;
assign img[ 4696] = 207;
assign img[ 4697] = 255;
assign img[ 4698] = 223;
assign img[ 4699] = 253;
assign img[ 4700] = 255;
assign img[ 4701] = 255;
assign img[ 4702] = 238;
assign img[ 4703] = 206;
assign img[ 4704] = 156;
assign img[ 4705] = 171;
assign img[ 4706] = 250;
assign img[ 4707] = 255;
assign img[ 4708] = 255;
assign img[ 4709] = 239;
assign img[ 4710] = 238;
assign img[ 4711] = 222;
assign img[ 4712] = 254;
assign img[ 4713] = 255;
assign img[ 4714] = 238;
assign img[ 4715] = 238;
assign img[ 4716] = 238;
assign img[ 4717] = 254;
assign img[ 4718] = 255;
assign img[ 4719] = 255;
assign img[ 4720] = 221;
assign img[ 4721] = 253;
assign img[ 4722] = 255;
assign img[ 4723] = 255;
assign img[ 4724] = 221;
assign img[ 4725] = 255;
assign img[ 4726] = 255;
assign img[ 4727] = 255;
assign img[ 4728] = 223;
assign img[ 4729] = 221;
assign img[ 4730] = 221;
assign img[ 4731] = 221;
assign img[ 4732] = 255;
assign img[ 4733] = 255;
assign img[ 4734] = 255;
assign img[ 4735] = 255;
assign img[ 4736] = 96;
assign img[ 4737] = 238;
assign img[ 4738] = 254;
assign img[ 4739] = 255;
assign img[ 4740] = 221;
assign img[ 4741] = 255;
assign img[ 4742] = 207;
assign img[ 4743] = 238;
assign img[ 4744] = 238;
assign img[ 4745] = 255;
assign img[ 4746] = 254;
assign img[ 4747] = 255;
assign img[ 4748] = 255;
assign img[ 4749] = 255;
assign img[ 4750] = 255;
assign img[ 4751] = 255;
assign img[ 4752] = 221;
assign img[ 4753] = 255;
assign img[ 4754] = 255;
assign img[ 4755] = 255;
assign img[ 4756] = 255;
assign img[ 4757] = 255;
assign img[ 4758] = 255;
assign img[ 4759] = 255;
assign img[ 4760] = 255;
assign img[ 4761] = 223;
assign img[ 4762] = 236;
assign img[ 4763] = 254;
assign img[ 4764] = 254;
assign img[ 4765] = 255;
assign img[ 4766] = 255;
assign img[ 4767] = 255;
assign img[ 4768] = 223;
assign img[ 4769] = 255;
assign img[ 4770] = 254;
assign img[ 4771] = 255;
assign img[ 4772] = 255;
assign img[ 4773] = 255;
assign img[ 4774] = 255;
assign img[ 4775] = 255;
assign img[ 4776] = 238;
assign img[ 4777] = 238;
assign img[ 4778] = 238;
assign img[ 4779] = 223;
assign img[ 4780] = 221;
assign img[ 4781] = 255;
assign img[ 4782] = 255;
assign img[ 4783] = 255;
assign img[ 4784] = 255;
assign img[ 4785] = 255;
assign img[ 4786] = 255;
assign img[ 4787] = 255;
assign img[ 4788] = 255;
assign img[ 4789] = 255;
assign img[ 4790] = 255;
assign img[ 4791] = 255;
assign img[ 4792] = 239;
assign img[ 4793] = 238;
assign img[ 4794] = 206;
assign img[ 4795] = 221;
assign img[ 4796] = 253;
assign img[ 4797] = 223;
assign img[ 4798] = 253;
assign img[ 4799] = 255;
assign img[ 4800] = 255;
assign img[ 4801] = 255;
assign img[ 4802] = 255;
assign img[ 4803] = 255;
assign img[ 4804] = 255;
assign img[ 4805] = 255;
assign img[ 4806] = 255;
assign img[ 4807] = 239;
assign img[ 4808] = 238;
assign img[ 4809] = 238;
assign img[ 4810] = 238;
assign img[ 4811] = 238;
assign img[ 4812] = 254;
assign img[ 4813] = 255;
assign img[ 4814] = 255;
assign img[ 4815] = 255;
assign img[ 4816] = 255;
assign img[ 4817] = 255;
assign img[ 4818] = 255;
assign img[ 4819] = 255;
assign img[ 4820] = 223;
assign img[ 4821] = 221;
assign img[ 4822] = 253;
assign img[ 4823] = 255;
assign img[ 4824] = 239;
assign img[ 4825] = 238;
assign img[ 4826] = 238;
assign img[ 4827] = 238;
assign img[ 4828] = 254;
assign img[ 4829] = 255;
assign img[ 4830] = 255;
assign img[ 4831] = 223;
assign img[ 4832] = 204;
assign img[ 4833] = 204;
assign img[ 4834] = 236;
assign img[ 4835] = 238;
assign img[ 4836] = 238;
assign img[ 4837] = 255;
assign img[ 4838] = 239;
assign img[ 4839] = 238;
assign img[ 4840] = 254;
assign img[ 4841] = 255;
assign img[ 4842] = 255;
assign img[ 4843] = 255;
assign img[ 4844] = 255;
assign img[ 4845] = 255;
assign img[ 4846] = 255;
assign img[ 4847] = 255;
assign img[ 4848] = 223;
assign img[ 4849] = 221;
assign img[ 4850] = 253;
assign img[ 4851] = 255;
assign img[ 4852] = 238;
assign img[ 4853] = 238;
assign img[ 4854] = 238;
assign img[ 4855] = 255;
assign img[ 4856] = 254;
assign img[ 4857] = 238;
assign img[ 4858] = 238;
assign img[ 4859] = 255;
assign img[ 4860] = 255;
assign img[ 4861] = 255;
assign img[ 4862] = 255;
assign img[ 4863] = 255;
assign img[ 4864] = 96;
assign img[ 4865] = 238;
assign img[ 4866] = 238;
assign img[ 4867] = 238;
assign img[ 4868] = 238;
assign img[ 4869] = 238;
assign img[ 4870] = 238;
assign img[ 4871] = 254;
assign img[ 4872] = 255;
assign img[ 4873] = 255;
assign img[ 4874] = 239;
assign img[ 4875] = 255;
assign img[ 4876] = 239;
assign img[ 4877] = 238;
assign img[ 4878] = 238;
assign img[ 4879] = 238;
assign img[ 4880] = 238;
assign img[ 4881] = 238;
assign img[ 4882] = 238;
assign img[ 4883] = 238;
assign img[ 4884] = 254;
assign img[ 4885] = 255;
assign img[ 4886] = 255;
assign img[ 4887] = 255;
assign img[ 4888] = 255;
assign img[ 4889] = 255;
assign img[ 4890] = 221;
assign img[ 4891] = 253;
assign img[ 4892] = 255;
assign img[ 4893] = 255;
assign img[ 4894] = 255;
assign img[ 4895] = 255;
assign img[ 4896] = 239;
assign img[ 4897] = 238;
assign img[ 4898] = 238;
assign img[ 4899] = 238;
assign img[ 4900] = 238;
assign img[ 4901] = 238;
assign img[ 4902] = 254;
assign img[ 4903] = 255;
assign img[ 4904] = 255;
assign img[ 4905] = 255;
assign img[ 4906] = 255;
assign img[ 4907] = 223;
assign img[ 4908] = 221;
assign img[ 4909] = 204;
assign img[ 4910] = 252;
assign img[ 4911] = 255;
assign img[ 4912] = 255;
assign img[ 4913] = 255;
assign img[ 4914] = 255;
assign img[ 4915] = 255;
assign img[ 4916] = 255;
assign img[ 4917] = 255;
assign img[ 4918] = 255;
assign img[ 4919] = 255;
assign img[ 4920] = 255;
assign img[ 4921] = 255;
assign img[ 4922] = 239;
assign img[ 4923] = 255;
assign img[ 4924] = 255;
assign img[ 4925] = 239;
assign img[ 4926] = 238;
assign img[ 4927] = 255;
assign img[ 4928] = 255;
assign img[ 4929] = 255;
assign img[ 4930] = 255;
assign img[ 4931] = 255;
assign img[ 4932] = 255;
assign img[ 4933] = 255;
assign img[ 4934] = 255;
assign img[ 4935] = 255;
assign img[ 4936] = 255;
assign img[ 4937] = 255;
assign img[ 4938] = 255;
assign img[ 4939] = 255;
assign img[ 4940] = 255;
assign img[ 4941] = 255;
assign img[ 4942] = 255;
assign img[ 4943] = 255;
assign img[ 4944] = 255;
assign img[ 4945] = 255;
assign img[ 4946] = 223;
assign img[ 4947] = 223;
assign img[ 4948] = 255;
assign img[ 4949] = 255;
assign img[ 4950] = 255;
assign img[ 4951] = 255;
assign img[ 4952] = 255;
assign img[ 4953] = 255;
assign img[ 4954] = 255;
assign img[ 4955] = 239;
assign img[ 4956] = 238;
assign img[ 4957] = 238;
assign img[ 4958] = 238;
assign img[ 4959] = 255;
assign img[ 4960] = 238;
assign img[ 4961] = 238;
assign img[ 4962] = 254;
assign img[ 4963] = 255;
assign img[ 4964] = 255;
assign img[ 4965] = 238;
assign img[ 4966] = 238;
assign img[ 4967] = 238;
assign img[ 4968] = 238;
assign img[ 4969] = 255;
assign img[ 4970] = 255;
assign img[ 4971] = 255;
assign img[ 4972] = 221;
assign img[ 4973] = 255;
assign img[ 4974] = 255;
assign img[ 4975] = 255;
assign img[ 4976] = 239;
assign img[ 4977] = 238;
assign img[ 4978] = 254;
assign img[ 4979] = 255;
assign img[ 4980] = 238;
assign img[ 4981] = 238;
assign img[ 4982] = 238;
assign img[ 4983] = 238;
assign img[ 4984] = 238;
assign img[ 4985] = 255;
assign img[ 4986] = 238;
assign img[ 4987] = 239;
assign img[ 4988] = 255;
assign img[ 4989] = 255;
assign img[ 4990] = 239;
assign img[ 4991] = 238;
assign img[ 4992] = 96;
assign img[ 4993] = 255;
assign img[ 4994] = 255;
assign img[ 4995] = 223;
assign img[ 4996] = 221;
assign img[ 4997] = 221;
assign img[ 4998] = 221;
assign img[ 4999] = 253;
assign img[ 5000] = 255;
assign img[ 5001] = 255;
assign img[ 5002] = 255;
assign img[ 5003] = 255;
assign img[ 5004] = 255;
assign img[ 5005] = 255;
assign img[ 5006] = 223;
assign img[ 5007] = 255;
assign img[ 5008] = 255;
assign img[ 5009] = 255;
assign img[ 5010] = 255;
assign img[ 5011] = 223;
assign img[ 5012] = 204;
assign img[ 5013] = 238;
assign img[ 5014] = 238;
assign img[ 5015] = 254;
assign img[ 5016] = 255;
assign img[ 5017] = 255;
assign img[ 5018] = 255;
assign img[ 5019] = 255;
assign img[ 5020] = 255;
assign img[ 5021] = 255;
assign img[ 5022] = 255;
assign img[ 5023] = 223;
assign img[ 5024] = 253;
assign img[ 5025] = 255;
assign img[ 5026] = 255;
assign img[ 5027] = 255;
assign img[ 5028] = 255;
assign img[ 5029] = 255;
assign img[ 5030] = 255;
assign img[ 5031] = 255;
assign img[ 5032] = 255;
assign img[ 5033] = 255;
assign img[ 5034] = 255;
assign img[ 5035] = 255;
assign img[ 5036] = 255;
assign img[ 5037] = 239;
assign img[ 5038] = 238;
assign img[ 5039] = 238;
assign img[ 5040] = 254;
assign img[ 5041] = 255;
assign img[ 5042] = 255;
assign img[ 5043] = 239;
assign img[ 5044] = 238;
assign img[ 5045] = 255;
assign img[ 5046] = 255;
assign img[ 5047] = 255;
assign img[ 5048] = 255;
assign img[ 5049] = 255;
assign img[ 5050] = 255;
assign img[ 5051] = 255;
assign img[ 5052] = 254;
assign img[ 5053] = 255;
assign img[ 5054] = 204;
assign img[ 5055] = 254;
assign img[ 5056] = 255;
assign img[ 5057] = 255;
assign img[ 5058] = 206;
assign img[ 5059] = 238;
assign img[ 5060] = 238;
assign img[ 5061] = 238;
assign img[ 5062] = 238;
assign img[ 5063] = 238;
assign img[ 5064] = 238;
assign img[ 5065] = 238;
assign img[ 5066] = 254;
assign img[ 5067] = 255;
assign img[ 5068] = 239;
assign img[ 5069] = 238;
assign img[ 5070] = 238;
assign img[ 5071] = 255;
assign img[ 5072] = 255;
assign img[ 5073] = 255;
assign img[ 5074] = 239;
assign img[ 5075] = 238;
assign img[ 5076] = 254;
assign img[ 5077] = 239;
assign img[ 5078] = 238;
assign img[ 5079] = 238;
assign img[ 5080] = 222;
assign img[ 5081] = 221;
assign img[ 5082] = 253;
assign img[ 5083] = 223;
assign img[ 5084] = 253;
assign img[ 5085] = 255;
assign img[ 5086] = 255;
assign img[ 5087] = 255;
assign img[ 5088] = 223;
assign img[ 5089] = 221;
assign img[ 5090] = 253;
assign img[ 5091] = 255;
assign img[ 5092] = 255;
assign img[ 5093] = 207;
assign img[ 5094] = 204;
assign img[ 5095] = 236;
assign img[ 5096] = 254;
assign img[ 5097] = 255;
assign img[ 5098] = 238;
assign img[ 5099] = 255;
assign img[ 5100] = 238;
assign img[ 5101] = 238;
assign img[ 5102] = 238;
assign img[ 5103] = 238;
assign img[ 5104] = 238;
assign img[ 5105] = 238;
assign img[ 5106] = 220;
assign img[ 5107] = 221;
assign img[ 5108] = 221;
assign img[ 5109] = 221;
assign img[ 5110] = 253;
assign img[ 5111] = 255;
assign img[ 5112] = 255;
assign img[ 5113] = 255;
assign img[ 5114] = 221;
assign img[ 5115] = 205;
assign img[ 5116] = 204;
assign img[ 5117] = 252;
assign img[ 5118] = 239;
assign img[ 5119] = 238;
assign img[ 5120] = 96;
assign img[ 5121] = 238;
assign img[ 5122] = 238;
assign img[ 5123] = 207;
assign img[ 5124] = 204;
assign img[ 5125] = 204;
assign img[ 5126] = 204;
assign img[ 5127] = 238;
assign img[ 5128] = 238;
assign img[ 5129] = 255;
assign img[ 5130] = 254;
assign img[ 5131] = 255;
assign img[ 5132] = 205;
assign img[ 5133] = 204;
assign img[ 5134] = 204;
assign img[ 5135] = 253;
assign img[ 5136] = 187;
assign img[ 5137] = 255;
assign img[ 5138] = 255;
assign img[ 5139] = 255;
assign img[ 5140] = 255;
assign img[ 5141] = 255;
assign img[ 5142] = 255;
assign img[ 5143] = 255;
assign img[ 5144] = 254;
assign img[ 5145] = 255;
assign img[ 5146] = 255;
assign img[ 5147] = 255;
assign img[ 5148] = 255;
assign img[ 5149] = 255;
assign img[ 5150] = 255;
assign img[ 5151] = 191;
assign img[ 5152] = 187;
assign img[ 5153] = 255;
assign img[ 5154] = 255;
assign img[ 5155] = 255;
assign img[ 5156] = 255;
assign img[ 5157] = 255;
assign img[ 5158] = 255;
assign img[ 5159] = 255;
assign img[ 5160] = 255;
assign img[ 5161] = 255;
assign img[ 5162] = 255;
assign img[ 5163] = 255;
assign img[ 5164] = 255;
assign img[ 5165] = 239;
assign img[ 5166] = 238;
assign img[ 5167] = 223;
assign img[ 5168] = 255;
assign img[ 5169] = 255;
assign img[ 5170] = 255;
assign img[ 5171] = 255;
assign img[ 5172] = 255;
assign img[ 5173] = 255;
assign img[ 5174] = 255;
assign img[ 5175] = 255;
assign img[ 5176] = 255;
assign img[ 5177] = 239;
assign img[ 5178] = 238;
assign img[ 5179] = 238;
assign img[ 5180] = 238;
assign img[ 5181] = 238;
assign img[ 5182] = 204;
assign img[ 5183] = 238;
assign img[ 5184] = 238;
assign img[ 5185] = 255;
assign img[ 5186] = 207;
assign img[ 5187] = 238;
assign img[ 5188] = 254;
assign img[ 5189] = 255;
assign img[ 5190] = 223;
assign img[ 5191] = 255;
assign img[ 5192] = 238;
assign img[ 5193] = 255;
assign img[ 5194] = 255;
assign img[ 5195] = 255;
assign img[ 5196] = 255;
assign img[ 5197] = 255;
assign img[ 5198] = 255;
assign img[ 5199] = 255;
assign img[ 5200] = 255;
assign img[ 5201] = 255;
assign img[ 5202] = 239;
assign img[ 5203] = 238;
assign img[ 5204] = 254;
assign img[ 5205] = 239;
assign img[ 5206] = 238;
assign img[ 5207] = 238;
assign img[ 5208] = 238;
assign img[ 5209] = 255;
assign img[ 5210] = 255;
assign img[ 5211] = 255;
assign img[ 5212] = 255;
assign img[ 5213] = 255;
assign img[ 5214] = 255;
assign img[ 5215] = 255;
assign img[ 5216] = 187;
assign img[ 5217] = 187;
assign img[ 5218] = 251;
assign img[ 5219] = 255;
assign img[ 5220] = 255;
assign img[ 5221] = 255;
assign img[ 5222] = 255;
assign img[ 5223] = 255;
assign img[ 5224] = 255;
assign img[ 5225] = 255;
assign img[ 5226] = 255;
assign img[ 5227] = 255;
assign img[ 5228] = 255;
assign img[ 5229] = 255;
assign img[ 5230] = 255;
assign img[ 5231] = 255;
assign img[ 5232] = 239;
assign img[ 5233] = 206;
assign img[ 5234] = 220;
assign img[ 5235] = 221;
assign img[ 5236] = 204;
assign img[ 5237] = 221;
assign img[ 5238] = 253;
assign img[ 5239] = 255;
assign img[ 5240] = 255;
assign img[ 5241] = 255;
assign img[ 5242] = 255;
assign img[ 5243] = 223;
assign img[ 5244] = 205;
assign img[ 5245] = 238;
assign img[ 5246] = 238;
assign img[ 5247] = 238;
assign img[ 5248] = 96;
assign img[ 5249] = 223;
assign img[ 5250] = 221;
assign img[ 5251] = 253;
assign img[ 5252] = 223;
assign img[ 5253] = 221;
assign img[ 5254] = 221;
assign img[ 5255] = 253;
assign img[ 5256] = 255;
assign img[ 5257] = 255;
assign img[ 5258] = 255;
assign img[ 5259] = 223;
assign img[ 5260] = 205;
assign img[ 5261] = 238;
assign img[ 5262] = 238;
assign img[ 5263] = 206;
assign img[ 5264] = 236;
assign img[ 5265] = 254;
assign img[ 5266] = 254;
assign img[ 5267] = 255;
assign img[ 5268] = 221;
assign img[ 5269] = 255;
assign img[ 5270] = 239;
assign img[ 5271] = 255;
assign img[ 5272] = 238;
assign img[ 5273] = 238;
assign img[ 5274] = 254;
assign img[ 5275] = 255;
assign img[ 5276] = 255;
assign img[ 5277] = 255;
assign img[ 5278] = 255;
assign img[ 5279] = 255;
assign img[ 5280] = 221;
assign img[ 5281] = 255;
assign img[ 5282] = 255;
assign img[ 5283] = 255;
assign img[ 5284] = 255;
assign img[ 5285] = 239;
assign img[ 5286] = 254;
assign img[ 5287] = 239;
assign img[ 5288] = 238;
assign img[ 5289] = 255;
assign img[ 5290] = 255;
assign img[ 5291] = 255;
assign img[ 5292] = 255;
assign img[ 5293] = 191;
assign img[ 5294] = 139;
assign img[ 5295] = 238;
assign img[ 5296] = 254;
assign img[ 5297] = 255;
assign img[ 5298] = 255;
assign img[ 5299] = 255;
assign img[ 5300] = 255;
assign img[ 5301] = 255;
assign img[ 5302] = 255;
assign img[ 5303] = 255;
assign img[ 5304] = 255;
assign img[ 5305] = 255;
assign img[ 5306] = 239;
assign img[ 5307] = 238;
assign img[ 5308] = 238;
assign img[ 5309] = 238;
assign img[ 5310] = 170;
assign img[ 5311] = 254;
assign img[ 5312] = 255;
assign img[ 5313] = 239;
assign img[ 5314] = 239;
assign img[ 5315] = 238;
assign img[ 5316] = 238;
assign img[ 5317] = 255;
assign img[ 5318] = 238;
assign img[ 5319] = 238;
assign img[ 5320] = 238;
assign img[ 5321] = 238;
assign img[ 5322] = 255;
assign img[ 5323] = 255;
assign img[ 5324] = 255;
assign img[ 5325] = 255;
assign img[ 5326] = 255;
assign img[ 5327] = 255;
assign img[ 5328] = 239;
assign img[ 5329] = 255;
assign img[ 5330] = 255;
assign img[ 5331] = 239;
assign img[ 5332] = 238;
assign img[ 5333] = 238;
assign img[ 5334] = 206;
assign img[ 5335] = 238;
assign img[ 5336] = 206;
assign img[ 5337] = 221;
assign img[ 5338] = 220;
assign img[ 5339] = 221;
assign img[ 5340] = 221;
assign img[ 5341] = 255;
assign img[ 5342] = 255;
assign img[ 5343] = 255;
assign img[ 5344] = 223;
assign img[ 5345] = 221;
assign img[ 5346] = 253;
assign img[ 5347] = 255;
assign img[ 5348] = 255;
assign img[ 5349] = 255;
assign img[ 5350] = 255;
assign img[ 5351] = 255;
assign img[ 5352] = 255;
assign img[ 5353] = 239;
assign img[ 5354] = 238;
assign img[ 5355] = 238;
assign img[ 5356] = 206;
assign img[ 5357] = 238;
assign img[ 5358] = 238;
assign img[ 5359] = 238;
assign img[ 5360] = 222;
assign img[ 5361] = 239;
assign img[ 5362] = 254;
assign img[ 5363] = 255;
assign img[ 5364] = 221;
assign img[ 5365] = 253;
assign img[ 5366] = 255;
assign img[ 5367] = 255;
assign img[ 5368] = 255;
assign img[ 5369] = 255;
assign img[ 5370] = 255;
assign img[ 5371] = 223;
assign img[ 5372] = 253;
assign img[ 5373] = 223;
assign img[ 5374] = 221;
assign img[ 5375] = 255;
assign img[ 5376] = 96;
assign img[ 5377] = 255;
assign img[ 5378] = 255;
assign img[ 5379] = 255;
assign img[ 5380] = 221;
assign img[ 5381] = 205;
assign img[ 5382] = 236;
assign img[ 5383] = 238;
assign img[ 5384] = 238;
assign img[ 5385] = 255;
assign img[ 5386] = 238;
assign img[ 5387] = 238;
assign img[ 5388] = 204;
assign img[ 5389] = 238;
assign img[ 5390] = 238;
assign img[ 5391] = 255;
assign img[ 5392] = 221;
assign img[ 5393] = 253;
assign img[ 5394] = 255;
assign img[ 5395] = 239;
assign img[ 5396] = 238;
assign img[ 5397] = 238;
assign img[ 5398] = 238;
assign img[ 5399] = 255;
assign img[ 5400] = 255;
assign img[ 5401] = 255;
assign img[ 5402] = 207;
assign img[ 5403] = 238;
assign img[ 5404] = 238;
assign img[ 5405] = 255;
assign img[ 5406] = 223;
assign img[ 5407] = 223;
assign img[ 5408] = 253;
assign img[ 5409] = 255;
assign img[ 5410] = 255;
assign img[ 5411] = 255;
assign img[ 5412] = 239;
assign img[ 5413] = 238;
assign img[ 5414] = 238;
assign img[ 5415] = 238;
assign img[ 5416] = 238;
assign img[ 5417] = 238;
assign img[ 5418] = 238;
assign img[ 5419] = 191;
assign img[ 5420] = 255;
assign img[ 5421] = 255;
assign img[ 5422] = 238;
assign img[ 5423] = 255;
assign img[ 5424] = 238;
assign img[ 5425] = 238;
assign img[ 5426] = 238;
assign img[ 5427] = 238;
assign img[ 5428] = 254;
assign img[ 5429] = 255;
assign img[ 5430] = 255;
assign img[ 5431] = 255;
assign img[ 5432] = 239;
assign img[ 5433] = 239;
assign img[ 5434] = 238;
assign img[ 5435] = 238;
assign img[ 5436] = 238;
assign img[ 5437] = 255;
assign img[ 5438] = 255;
assign img[ 5439] = 255;
assign img[ 5440] = 255;
assign img[ 5441] = 255;
assign img[ 5442] = 255;
assign img[ 5443] = 255;
assign img[ 5444] = 255;
assign img[ 5445] = 255;
assign img[ 5446] = 255;
assign img[ 5447] = 239;
assign img[ 5448] = 238;
assign img[ 5449] = 238;
assign img[ 5450] = 254;
assign img[ 5451] = 255;
assign img[ 5452] = 255;
assign img[ 5453] = 255;
assign img[ 5454] = 238;
assign img[ 5455] = 254;
assign img[ 5456] = 238;
assign img[ 5457] = 238;
assign img[ 5458] = 238;
assign img[ 5459] = 238;
assign img[ 5460] = 174;
assign img[ 5461] = 255;
assign img[ 5462] = 255;
assign img[ 5463] = 255;
assign img[ 5464] = 255;
assign img[ 5465] = 255;
assign img[ 5466] = 255;
assign img[ 5467] = 255;
assign img[ 5468] = 238;
assign img[ 5469] = 238;
assign img[ 5470] = 255;
assign img[ 5471] = 207;
assign img[ 5472] = 220;
assign img[ 5473] = 221;
assign img[ 5474] = 253;
assign img[ 5475] = 255;
assign img[ 5476] = 255;
assign img[ 5477] = 223;
assign img[ 5478] = 204;
assign img[ 5479] = 236;
assign img[ 5480] = 238;
assign img[ 5481] = 238;
assign img[ 5482] = 238;
assign img[ 5483] = 255;
assign img[ 5484] = 255;
assign img[ 5485] = 255;
assign img[ 5486] = 255;
assign img[ 5487] = 255;
assign img[ 5488] = 255;
assign img[ 5489] = 255;
assign img[ 5490] = 255;
assign img[ 5491] = 255;
assign img[ 5492] = 223;
assign img[ 5493] = 223;
assign img[ 5494] = 255;
assign img[ 5495] = 255;
assign img[ 5496] = 255;
assign img[ 5497] = 255;
assign img[ 5498] = 155;
assign img[ 5499] = 223;
assign img[ 5500] = 238;
assign img[ 5501] = 255;
assign img[ 5502] = 239;
assign img[ 5503] = 238;
assign img[ 5504] = 96;
assign img[ 5505] = 255;
assign img[ 5506] = 255;
assign img[ 5507] = 255;
assign img[ 5508] = 255;
assign img[ 5509] = 239;
assign img[ 5510] = 239;
assign img[ 5511] = 238;
assign img[ 5512] = 238;
assign img[ 5513] = 254;
assign img[ 5514] = 255;
assign img[ 5515] = 206;
assign img[ 5516] = 204;
assign img[ 5517] = 220;
assign img[ 5518] = 221;
assign img[ 5519] = 255;
assign img[ 5520] = 255;
assign img[ 5521] = 255;
assign img[ 5522] = 255;
assign img[ 5523] = 223;
assign img[ 5524] = 236;
assign img[ 5525] = 238;
assign img[ 5526] = 238;
assign img[ 5527] = 255;
assign img[ 5528] = 255;
assign img[ 5529] = 255;
assign img[ 5530] = 239;
assign img[ 5531] = 238;
assign img[ 5532] = 238;
assign img[ 5533] = 238;
assign img[ 5534] = 238;
assign img[ 5535] = 174;
assign img[ 5536] = 136;
assign img[ 5537] = 255;
assign img[ 5538] = 255;
assign img[ 5539] = 255;
assign img[ 5540] = 223;
assign img[ 5541] = 255;
assign img[ 5542] = 254;
assign img[ 5543] = 238;
assign img[ 5544] = 238;
assign img[ 5545] = 238;
assign img[ 5546] = 238;
assign img[ 5547] = 254;
assign img[ 5548] = 255;
assign img[ 5549] = 239;
assign img[ 5550] = 238;
assign img[ 5551] = 223;
assign img[ 5552] = 255;
assign img[ 5553] = 255;
assign img[ 5554] = 239;
assign img[ 5555] = 206;
assign img[ 5556] = 254;
assign img[ 5557] = 255;
assign img[ 5558] = 207;
assign img[ 5559] = 238;
assign img[ 5560] = 254;
assign img[ 5561] = 255;
assign img[ 5562] = 255;
assign img[ 5563] = 255;
assign img[ 5564] = 255;
assign img[ 5565] = 239;
assign img[ 5566] = 238;
assign img[ 5567] = 255;
assign img[ 5568] = 255;
assign img[ 5569] = 255;
assign img[ 5570] = 255;
assign img[ 5571] = 255;
assign img[ 5572] = 255;
assign img[ 5573] = 255;
assign img[ 5574] = 238;
assign img[ 5575] = 255;
assign img[ 5576] = 255;
assign img[ 5577] = 239;
assign img[ 5578] = 254;
assign img[ 5579] = 255;
assign img[ 5580] = 223;
assign img[ 5581] = 221;
assign img[ 5582] = 236;
assign img[ 5583] = 254;
assign img[ 5584] = 206;
assign img[ 5585] = 255;
assign img[ 5586] = 238;
assign img[ 5587] = 255;
assign img[ 5588] = 254;
assign img[ 5589] = 255;
assign img[ 5590] = 238;
assign img[ 5591] = 238;
assign img[ 5592] = 238;
assign img[ 5593] = 238;
assign img[ 5594] = 255;
assign img[ 5595] = 255;
assign img[ 5596] = 255;
assign img[ 5597] = 255;
assign img[ 5598] = 255;
assign img[ 5599] = 255;
assign img[ 5600] = 155;
assign img[ 5601] = 153;
assign img[ 5602] = 232;
assign img[ 5603] = 254;
assign img[ 5604] = 255;
assign img[ 5605] = 255;
assign img[ 5606] = 238;
assign img[ 5607] = 238;
assign img[ 5608] = 238;
assign img[ 5609] = 254;
assign img[ 5610] = 238;
assign img[ 5611] = 255;
assign img[ 5612] = 206;
assign img[ 5613] = 254;
assign img[ 5614] = 255;
assign img[ 5615] = 255;
assign img[ 5616] = 223;
assign img[ 5617] = 221;
assign img[ 5618] = 253;
assign img[ 5619] = 255;
assign img[ 5620] = 255;
assign img[ 5621] = 239;
assign img[ 5622] = 238;
assign img[ 5623] = 238;
assign img[ 5624] = 254;
assign img[ 5625] = 239;
assign img[ 5626] = 170;
assign img[ 5627] = 206;
assign img[ 5628] = 220;
assign img[ 5629] = 255;
assign img[ 5630] = 255;
assign img[ 5631] = 255;
assign img[ 5632] = 96;
assign img[ 5633] = 238;
assign img[ 5634] = 254;
assign img[ 5635] = 239;
assign img[ 5636] = 238;
assign img[ 5637] = 238;
assign img[ 5638] = 254;
assign img[ 5639] = 255;
assign img[ 5640] = 255;
assign img[ 5641] = 254;
assign img[ 5642] = 254;
assign img[ 5643] = 255;
assign img[ 5644] = 255;
assign img[ 5645] = 255;
assign img[ 5646] = 223;
assign img[ 5647] = 239;
assign img[ 5648] = 222;
assign img[ 5649] = 205;
assign img[ 5650] = 236;
assign img[ 5651] = 206;
assign img[ 5652] = 204;
assign img[ 5653] = 238;
assign img[ 5654] = 238;
assign img[ 5655] = 238;
assign img[ 5656] = 255;
assign img[ 5657] = 191;
assign img[ 5658] = 223;
assign img[ 5659] = 255;
assign img[ 5660] = 255;
assign img[ 5661] = 255;
assign img[ 5662] = 255;
assign img[ 5663] = 255;
assign img[ 5664] = 255;
assign img[ 5665] = 255;
assign img[ 5666] = 255;
assign img[ 5667] = 255;
assign img[ 5668] = 255;
assign img[ 5669] = 255;
assign img[ 5670] = 255;
assign img[ 5671] = 255;
assign img[ 5672] = 255;
assign img[ 5673] = 255;
assign img[ 5674] = 239;
assign img[ 5675] = 238;
assign img[ 5676] = 238;
assign img[ 5677] = 238;
assign img[ 5678] = 238;
assign img[ 5679] = 238;
assign img[ 5680] = 238;
assign img[ 5681] = 255;
assign img[ 5682] = 238;
assign img[ 5683] = 254;
assign img[ 5684] = 255;
assign img[ 5685] = 255;
assign img[ 5686] = 255;
assign img[ 5687] = 255;
assign img[ 5688] = 239;
assign img[ 5689] = 238;
assign img[ 5690] = 238;
assign img[ 5691] = 254;
assign img[ 5692] = 255;
assign img[ 5693] = 223;
assign img[ 5694] = 238;
assign img[ 5695] = 255;
assign img[ 5696] = 255;
assign img[ 5697] = 255;
assign img[ 5698] = 223;
assign img[ 5699] = 255;
assign img[ 5700] = 255;
assign img[ 5701] = 239;
assign img[ 5702] = 238;
assign img[ 5703] = 239;
assign img[ 5704] = 238;
assign img[ 5705] = 238;
assign img[ 5706] = 254;
assign img[ 5707] = 255;
assign img[ 5708] = 255;
assign img[ 5709] = 255;
assign img[ 5710] = 238;
assign img[ 5711] = 238;
assign img[ 5712] = 238;
assign img[ 5713] = 238;
assign img[ 5714] = 238;
assign img[ 5715] = 254;
assign img[ 5716] = 238;
assign img[ 5717] = 238;
assign img[ 5718] = 238;
assign img[ 5719] = 239;
assign img[ 5720] = 238;
assign img[ 5721] = 254;
assign img[ 5722] = 255;
assign img[ 5723] = 255;
assign img[ 5724] = 255;
assign img[ 5725] = 255;
assign img[ 5726] = 255;
assign img[ 5727] = 223;
assign img[ 5728] = 253;
assign img[ 5729] = 255;
assign img[ 5730] = 255;
assign img[ 5731] = 255;
assign img[ 5732] = 255;
assign img[ 5733] = 255;
assign img[ 5734] = 255;
assign img[ 5735] = 255;
assign img[ 5736] = 255;
assign img[ 5737] = 255;
assign img[ 5738] = 255;
assign img[ 5739] = 255;
assign img[ 5740] = 223;
assign img[ 5741] = 255;
assign img[ 5742] = 255;
assign img[ 5743] = 223;
assign img[ 5744] = 221;
assign img[ 5745] = 205;
assign img[ 5746] = 238;
assign img[ 5747] = 238;
assign img[ 5748] = 238;
assign img[ 5749] = 238;
assign img[ 5750] = 254;
assign img[ 5751] = 255;
assign img[ 5752] = 255;
assign img[ 5753] = 255;
assign img[ 5754] = 255;
assign img[ 5755] = 255;
assign img[ 5756] = 255;
assign img[ 5757] = 255;
assign img[ 5758] = 255;
assign img[ 5759] = 255;
assign img[ 5760] = 96;
assign img[ 5761] = 255;
assign img[ 5762] = 255;
assign img[ 5763] = 255;
assign img[ 5764] = 255;
assign img[ 5765] = 207;
assign img[ 5766] = 204;
assign img[ 5767] = 238;
assign img[ 5768] = 238;
assign img[ 5769] = 238;
assign img[ 5770] = 238;
assign img[ 5771] = 238;
assign img[ 5772] = 238;
assign img[ 5773] = 238;
assign img[ 5774] = 204;
assign img[ 5775] = 236;
assign img[ 5776] = 254;
assign img[ 5777] = 255;
assign img[ 5778] = 255;
assign img[ 5779] = 255;
assign img[ 5780] = 238;
assign img[ 5781] = 254;
assign img[ 5782] = 206;
assign img[ 5783] = 255;
assign img[ 5784] = 254;
assign img[ 5785] = 190;
assign img[ 5786] = 187;
assign img[ 5787] = 255;
assign img[ 5788] = 254;
assign img[ 5789] = 255;
assign img[ 5790] = 239;
assign img[ 5791] = 174;
assign img[ 5792] = 238;
assign img[ 5793] = 238;
assign img[ 5794] = 238;
assign img[ 5795] = 255;
assign img[ 5796] = 255;
assign img[ 5797] = 255;
assign img[ 5798] = 255;
assign img[ 5799] = 239;
assign img[ 5800] = 238;
assign img[ 5801] = 238;
assign img[ 5802] = 206;
assign img[ 5803] = 174;
assign img[ 5804] = 238;
assign img[ 5805] = 255;
assign img[ 5806] = 255;
assign img[ 5807] = 255;
assign img[ 5808] = 255;
assign img[ 5809] = 255;
assign img[ 5810] = 255;
assign img[ 5811] = 255;
assign img[ 5812] = 255;
assign img[ 5813] = 255;
assign img[ 5814] = 255;
assign img[ 5815] = 255;
assign img[ 5816] = 255;
assign img[ 5817] = 255;
assign img[ 5818] = 255;
assign img[ 5819] = 255;
assign img[ 5820] = 255;
assign img[ 5821] = 255;
assign img[ 5822] = 255;
assign img[ 5823] = 255;
assign img[ 5824] = 255;
assign img[ 5825] = 255;
assign img[ 5826] = 255;
assign img[ 5827] = 255;
assign img[ 5828] = 255;
assign img[ 5829] = 255;
assign img[ 5830] = 255;
assign img[ 5831] = 239;
assign img[ 5832] = 238;
assign img[ 5833] = 238;
assign img[ 5834] = 254;
assign img[ 5835] = 255;
assign img[ 5836] = 255;
assign img[ 5837] = 255;
assign img[ 5838] = 255;
assign img[ 5839] = 255;
assign img[ 5840] = 239;
assign img[ 5841] = 238;
assign img[ 5842] = 238;
assign img[ 5843] = 238;
assign img[ 5844] = 174;
assign img[ 5845] = 138;
assign img[ 5846] = 234;
assign img[ 5847] = 238;
assign img[ 5848] = 206;
assign img[ 5849] = 221;
assign img[ 5850] = 253;
assign img[ 5851] = 255;
assign img[ 5852] = 255;
assign img[ 5853] = 255;
assign img[ 5854] = 255;
assign img[ 5855] = 207;
assign img[ 5856] = 236;
assign img[ 5857] = 239;
assign img[ 5858] = 255;
assign img[ 5859] = 255;
assign img[ 5860] = 255;
assign img[ 5861] = 239;
assign img[ 5862] = 254;
assign img[ 5863] = 255;
assign img[ 5864] = 255;
assign img[ 5865] = 255;
assign img[ 5866] = 255;
assign img[ 5867] = 255;
assign img[ 5868] = 255;
assign img[ 5869] = 255;
assign img[ 5870] = 255;
assign img[ 5871] = 239;
assign img[ 5872] = 238;
assign img[ 5873] = 206;
assign img[ 5874] = 220;
assign img[ 5875] = 239;
assign img[ 5876] = 254;
assign img[ 5877] = 255;
assign img[ 5878] = 255;
assign img[ 5879] = 255;
assign img[ 5880] = 255;
assign img[ 5881] = 255;
assign img[ 5882] = 255;
assign img[ 5883] = 255;
assign img[ 5884] = 255;
assign img[ 5885] = 255;
assign img[ 5886] = 239;
assign img[ 5887] = 238;
assign img[ 5888] = 96;
assign img[ 5889] = 238;
assign img[ 5890] = 254;
assign img[ 5891] = 255;
assign img[ 5892] = 239;
assign img[ 5893] = 238;
assign img[ 5894] = 206;
assign img[ 5895] = 238;
assign img[ 5896] = 238;
assign img[ 5897] = 255;
assign img[ 5898] = 255;
assign img[ 5899] = 255;
assign img[ 5900] = 255;
assign img[ 5901] = 255;
assign img[ 5902] = 255;
assign img[ 5903] = 255;
assign img[ 5904] = 238;
assign img[ 5905] = 238;
assign img[ 5906] = 254;
assign img[ 5907] = 223;
assign img[ 5908] = 221;
assign img[ 5909] = 253;
assign img[ 5910] = 206;
assign img[ 5911] = 238;
assign img[ 5912] = 254;
assign img[ 5913] = 221;
assign img[ 5914] = 221;
assign img[ 5915] = 253;
assign img[ 5916] = 255;
assign img[ 5917] = 255;
assign img[ 5918] = 239;
assign img[ 5919] = 238;
assign img[ 5920] = 186;
assign img[ 5921] = 255;
assign img[ 5922] = 255;
assign img[ 5923] = 255;
assign img[ 5924] = 255;
assign img[ 5925] = 255;
assign img[ 5926] = 255;
assign img[ 5927] = 255;
assign img[ 5928] = 255;
assign img[ 5929] = 255;
assign img[ 5930] = 255;
assign img[ 5931] = 255;
assign img[ 5932] = 205;
assign img[ 5933] = 238;
assign img[ 5934] = 238;
assign img[ 5935] = 238;
assign img[ 5936] = 254;
assign img[ 5937] = 255;
assign img[ 5938] = 255;
assign img[ 5939] = 255;
assign img[ 5940] = 255;
assign img[ 5941] = 255;
assign img[ 5942] = 255;
assign img[ 5943] = 255;
assign img[ 5944] = 255;
assign img[ 5945] = 255;
assign img[ 5946] = 255;
assign img[ 5947] = 255;
assign img[ 5948] = 238;
assign img[ 5949] = 238;
assign img[ 5950] = 254;
assign img[ 5951] = 255;
assign img[ 5952] = 255;
assign img[ 5953] = 255;
assign img[ 5954] = 255;
assign img[ 5955] = 255;
assign img[ 5956] = 255;
assign img[ 5957] = 255;
assign img[ 5958] = 255;
assign img[ 5959] = 255;
assign img[ 5960] = 255;
assign img[ 5961] = 255;
assign img[ 5962] = 255;
assign img[ 5963] = 255;
assign img[ 5964] = 255;
assign img[ 5965] = 255;
assign img[ 5966] = 255;
assign img[ 5967] = 255;
assign img[ 5968] = 255;
assign img[ 5969] = 255;
assign img[ 5970] = 223;
assign img[ 5971] = 204;
assign img[ 5972] = 204;
assign img[ 5973] = 221;
assign img[ 5974] = 253;
assign img[ 5975] = 255;
assign img[ 5976] = 255;
assign img[ 5977] = 255;
assign img[ 5978] = 255;
assign img[ 5979] = 239;
assign img[ 5980] = 238;
assign img[ 5981] = 238;
assign img[ 5982] = 238;
assign img[ 5983] = 206;
assign img[ 5984] = 238;
assign img[ 5985] = 255;
assign img[ 5986] = 255;
assign img[ 5987] = 255;
assign img[ 5988] = 255;
assign img[ 5989] = 239;
assign img[ 5990] = 238;
assign img[ 5991] = 206;
assign img[ 5992] = 236;
assign img[ 5993] = 255;
assign img[ 5994] = 255;
assign img[ 5995] = 223;
assign img[ 5996] = 221;
assign img[ 5997] = 253;
assign img[ 5998] = 255;
assign img[ 5999] = 255;
assign img[ 6000] = 239;
assign img[ 6001] = 238;
assign img[ 6002] = 238;
assign img[ 6003] = 238;
assign img[ 6004] = 238;
assign img[ 6005] = 238;
assign img[ 6006] = 204;
assign img[ 6007] = 254;
assign img[ 6008] = 238;
assign img[ 6009] = 255;
assign img[ 6010] = 255;
assign img[ 6011] = 223;
assign img[ 6012] = 221;
assign img[ 6013] = 253;
assign img[ 6014] = 255;
assign img[ 6015] = 255;
assign img[ 6016] = 96;
assign img[ 6017] = 223;
assign img[ 6018] = 253;
assign img[ 6019] = 255;
assign img[ 6020] = 255;
assign img[ 6021] = 255;
assign img[ 6022] = 255;
assign img[ 6023] = 255;
assign img[ 6024] = 255;
assign img[ 6025] = 255;
assign img[ 6026] = 255;
assign img[ 6027] = 255;
assign img[ 6028] = 255;
assign img[ 6029] = 255;
assign img[ 6030] = 159;
assign img[ 6031] = 171;
assign img[ 6032] = 234;
assign img[ 6033] = 255;
assign img[ 6034] = 255;
assign img[ 6035] = 255;
assign img[ 6036] = 187;
assign img[ 6037] = 255;
assign img[ 6038] = 255;
assign img[ 6039] = 255;
assign img[ 6040] = 255;
assign img[ 6041] = 239;
assign img[ 6042] = 204;
assign img[ 6043] = 254;
assign img[ 6044] = 254;
assign img[ 6045] = 254;
assign img[ 6046] = 238;
assign img[ 6047] = 238;
assign img[ 6048] = 170;
assign img[ 6049] = 255;
assign img[ 6050] = 255;
assign img[ 6051] = 255;
assign img[ 6052] = 255;
assign img[ 6053] = 255;
assign img[ 6054] = 255;
assign img[ 6055] = 255;
assign img[ 6056] = 255;
assign img[ 6057] = 255;
assign img[ 6058] = 239;
assign img[ 6059] = 238;
assign img[ 6060] = 255;
assign img[ 6061] = 239;
assign img[ 6062] = 238;
assign img[ 6063] = 255;
assign img[ 6064] = 255;
assign img[ 6065] = 255;
assign img[ 6066] = 255;
assign img[ 6067] = 255;
assign img[ 6068] = 255;
assign img[ 6069] = 255;
assign img[ 6070] = 255;
assign img[ 6071] = 255;
assign img[ 6072] = 255;
assign img[ 6073] = 255;
assign img[ 6074] = 255;
assign img[ 6075] = 255;
assign img[ 6076] = 255;
assign img[ 6077] = 255;
assign img[ 6078] = 255;
assign img[ 6079] = 255;
assign img[ 6080] = 255;
assign img[ 6081] = 255;
assign img[ 6082] = 255;
assign img[ 6083] = 255;
assign img[ 6084] = 255;
assign img[ 6085] = 239;
assign img[ 6086] = 238;
assign img[ 6087] = 238;
assign img[ 6088] = 238;
assign img[ 6089] = 238;
assign img[ 6090] = 238;
assign img[ 6091] = 238;
assign img[ 6092] = 254;
assign img[ 6093] = 255;
assign img[ 6094] = 255;
assign img[ 6095] = 255;
assign img[ 6096] = 255;
assign img[ 6097] = 255;
assign img[ 6098] = 255;
assign img[ 6099] = 255;
assign img[ 6100] = 207;
assign img[ 6101] = 204;
assign img[ 6102] = 236;
assign img[ 6103] = 238;
assign img[ 6104] = 238;
assign img[ 6105] = 238;
assign img[ 6106] = 223;
assign img[ 6107] = 221;
assign img[ 6108] = 253;
assign img[ 6109] = 255;
assign img[ 6110] = 255;
assign img[ 6111] = 255;
assign img[ 6112] = 255;
assign img[ 6113] = 239;
assign img[ 6114] = 238;
assign img[ 6115] = 238;
assign img[ 6116] = 238;
assign img[ 6117] = 238;
assign img[ 6118] = 238;
assign img[ 6119] = 238;
assign img[ 6120] = 254;
assign img[ 6121] = 255;
assign img[ 6122] = 238;
assign img[ 6123] = 238;
assign img[ 6124] = 238;
assign img[ 6125] = 238;
assign img[ 6126] = 238;
assign img[ 6127] = 254;
assign img[ 6128] = 255;
assign img[ 6129] = 159;
assign img[ 6130] = 221;
assign img[ 6131] = 255;
assign img[ 6132] = 255;
assign img[ 6133] = 255;
assign img[ 6134] = 238;
assign img[ 6135] = 238;
assign img[ 6136] = 238;
assign img[ 6137] = 255;
assign img[ 6138] = 255;
assign img[ 6139] = 255;
assign img[ 6140] = 255;
assign img[ 6141] = 255;
assign img[ 6142] = 223;
assign img[ 6143] = 255;
assign img[ 6144] = 96;
assign img[ 6145] = 206;
assign img[ 6146] = 236;
assign img[ 6147] = 206;
assign img[ 6148] = 252;
assign img[ 6149] = 254;
assign img[ 6150] = 255;
assign img[ 6151] = 255;
assign img[ 6152] = 255;
assign img[ 6153] = 255;
assign img[ 6154] = 255;
assign img[ 6155] = 191;
assign img[ 6156] = 186;
assign img[ 6157] = 255;
assign img[ 6158] = 254;
assign img[ 6159] = 255;
assign img[ 6160] = 206;
assign img[ 6161] = 204;
assign img[ 6162] = 252;
assign img[ 6163] = 223;
assign img[ 6164] = 236;
assign img[ 6165] = 238;
assign img[ 6166] = 238;
assign img[ 6167] = 254;
assign img[ 6168] = 254;
assign img[ 6169] = 238;
assign img[ 6170] = 238;
assign img[ 6171] = 238;
assign img[ 6172] = 238;
assign img[ 6173] = 255;
assign img[ 6174] = 223;
assign img[ 6175] = 221;
assign img[ 6176] = 237;
assign img[ 6177] = 238;
assign img[ 6178] = 254;
assign img[ 6179] = 255;
assign img[ 6180] = 255;
assign img[ 6181] = 255;
assign img[ 6182] = 255;
assign img[ 6183] = 255;
assign img[ 6184] = 238;
assign img[ 6185] = 238;
assign img[ 6186] = 206;
assign img[ 6187] = 238;
assign img[ 6188] = 238;
assign img[ 6189] = 255;
assign img[ 6190] = 255;
assign img[ 6191] = 223;
assign img[ 6192] = 255;
assign img[ 6193] = 239;
assign img[ 6194] = 206;
assign img[ 6195] = 238;
assign img[ 6196] = 254;
assign img[ 6197] = 255;
assign img[ 6198] = 255;
assign img[ 6199] = 255;
assign img[ 6200] = 253;
assign img[ 6201] = 255;
assign img[ 6202] = 221;
assign img[ 6203] = 255;
assign img[ 6204] = 255;
assign img[ 6205] = 255;
assign img[ 6206] = 255;
assign img[ 6207] = 255;
assign img[ 6208] = 255;
assign img[ 6209] = 255;
assign img[ 6210] = 255;
assign img[ 6211] = 255;
assign img[ 6212] = 255;
assign img[ 6213] = 255;
assign img[ 6214] = 239;
assign img[ 6215] = 255;
assign img[ 6216] = 255;
assign img[ 6217] = 255;
assign img[ 6218] = 255;
assign img[ 6219] = 255;
assign img[ 6220] = 255;
assign img[ 6221] = 255;
assign img[ 6222] = 221;
assign img[ 6223] = 255;
assign img[ 6224] = 255;
assign img[ 6225] = 255;
assign img[ 6226] = 255;
assign img[ 6227] = 255;
assign img[ 6228] = 255;
assign img[ 6229] = 223;
assign img[ 6230] = 238;
assign img[ 6231] = 238;
assign img[ 6232] = 238;
assign img[ 6233] = 254;
assign img[ 6234] = 255;
assign img[ 6235] = 255;
assign img[ 6236] = 255;
assign img[ 6237] = 255;
assign img[ 6238] = 255;
assign img[ 6239] = 255;
assign img[ 6240] = 255;
assign img[ 6241] = 223;
assign img[ 6242] = 253;
assign img[ 6243] = 255;
assign img[ 6244] = 255;
assign img[ 6245] = 239;
assign img[ 6246] = 206;
assign img[ 6247] = 254;
assign img[ 6248] = 238;
assign img[ 6249] = 238;
assign img[ 6250] = 238;
assign img[ 6251] = 238;
assign img[ 6252] = 206;
assign img[ 6253] = 254;
assign img[ 6254] = 255;
assign img[ 6255] = 255;
assign img[ 6256] = 238;
assign img[ 6257] = 238;
assign img[ 6258] = 238;
assign img[ 6259] = 255;
assign img[ 6260] = 191;
assign img[ 6261] = 187;
assign img[ 6262] = 217;
assign img[ 6263] = 255;
assign img[ 6264] = 255;
assign img[ 6265] = 255;
assign img[ 6266] = 255;
assign img[ 6267] = 239;
assign img[ 6268] = 206;
assign img[ 6269] = 238;
assign img[ 6270] = 206;
assign img[ 6271] = 236;
assign img[ 6272] = 96;
assign img[ 6273] = 206;
assign img[ 6274] = 252;
assign img[ 6275] = 255;
assign img[ 6276] = 255;
assign img[ 6277] = 255;
assign img[ 6278] = 207;
assign img[ 6279] = 238;
assign img[ 6280] = 238;
assign img[ 6281] = 238;
assign img[ 6282] = 238;
assign img[ 6283] = 238;
assign img[ 6284] = 238;
assign img[ 6285] = 238;
assign img[ 6286] = 206;
assign img[ 6287] = 204;
assign img[ 6288] = 252;
assign img[ 6289] = 255;
assign img[ 6290] = 255;
assign img[ 6291] = 255;
assign img[ 6292] = 223;
assign img[ 6293] = 255;
assign img[ 6294] = 223;
assign img[ 6295] = 253;
assign img[ 6296] = 255;
assign img[ 6297] = 255;
assign img[ 6298] = 255;
assign img[ 6299] = 255;
assign img[ 6300] = 255;
assign img[ 6301] = 255;
assign img[ 6302] = 255;
assign img[ 6303] = 255;
assign img[ 6304] = 155;
assign img[ 6305] = 171;
assign img[ 6306] = 238;
assign img[ 6307] = 255;
assign img[ 6308] = 223;
assign img[ 6309] = 255;
assign img[ 6310] = 255;
assign img[ 6311] = 255;
assign img[ 6312] = 238;
assign img[ 6313] = 238;
assign img[ 6314] = 222;
assign img[ 6315] = 255;
assign img[ 6316] = 255;
assign img[ 6317] = 223;
assign img[ 6318] = 253;
assign img[ 6319] = 255;
assign img[ 6320] = 255;
assign img[ 6321] = 223;
assign img[ 6322] = 221;
assign img[ 6323] = 255;
assign img[ 6324] = 255;
assign img[ 6325] = 255;
assign img[ 6326] = 255;
assign img[ 6327] = 255;
assign img[ 6328] = 255;
assign img[ 6329] = 239;
assign img[ 6330] = 206;
assign img[ 6331] = 204;
assign img[ 6332] = 252;
assign img[ 6333] = 255;
assign img[ 6334] = 255;
assign img[ 6335] = 255;
assign img[ 6336] = 255;
assign img[ 6337] = 255;
assign img[ 6338] = 255;
assign img[ 6339] = 255;
assign img[ 6340] = 207;
assign img[ 6341] = 204;
assign img[ 6342] = 204;
assign img[ 6343] = 238;
assign img[ 6344] = 238;
assign img[ 6345] = 238;
assign img[ 6346] = 238;
assign img[ 6347] = 238;
assign img[ 6348] = 238;
assign img[ 6349] = 239;
assign img[ 6350] = 255;
assign img[ 6351] = 255;
assign img[ 6352] = 239;
assign img[ 6353] = 238;
assign img[ 6354] = 238;
assign img[ 6355] = 238;
assign img[ 6356] = 238;
assign img[ 6357] = 206;
assign img[ 6358] = 238;
assign img[ 6359] = 238;
assign img[ 6360] = 238;
assign img[ 6361] = 238;
assign img[ 6362] = 238;
assign img[ 6363] = 255;
assign img[ 6364] = 255;
assign img[ 6365] = 255;
assign img[ 6366] = 255;
assign img[ 6367] = 239;
assign img[ 6368] = 204;
assign img[ 6369] = 238;
assign img[ 6370] = 254;
assign img[ 6371] = 239;
assign img[ 6372] = 238;
assign img[ 6373] = 255;
assign img[ 6374] = 191;
assign img[ 6375] = 255;
assign img[ 6376] = 255;
assign img[ 6377] = 255;
assign img[ 6378] = 255;
assign img[ 6379] = 223;
assign img[ 6380] = 255;
assign img[ 6381] = 255;
assign img[ 6382] = 255;
assign img[ 6383] = 255;
assign img[ 6384] = 223;
assign img[ 6385] = 221;
assign img[ 6386] = 253;
assign img[ 6387] = 255;
assign img[ 6388] = 255;
assign img[ 6389] = 239;
assign img[ 6390] = 238;
assign img[ 6391] = 238;
assign img[ 6392] = 238;
assign img[ 6393] = 255;
assign img[ 6394] = 238;
assign img[ 6395] = 238;
assign img[ 6396] = 254;
assign img[ 6397] = 255;
assign img[ 6398] = 223;
assign img[ 6399] = 255;
assign img[ 6400] = 96;
assign img[ 6401] = 238;
assign img[ 6402] = 238;
assign img[ 6403] = 255;
assign img[ 6404] = 239;
assign img[ 6405] = 238;
assign img[ 6406] = 254;
assign img[ 6407] = 255;
assign img[ 6408] = 239;
assign img[ 6409] = 255;
assign img[ 6410] = 254;
assign img[ 6411] = 255;
assign img[ 6412] = 221;
assign img[ 6413] = 255;
assign img[ 6414] = 255;
assign img[ 6415] = 255;
assign img[ 6416] = 238;
assign img[ 6417] = 254;
assign img[ 6418] = 255;
assign img[ 6419] = 255;
assign img[ 6420] = 238;
assign img[ 6421] = 238;
assign img[ 6422] = 254;
assign img[ 6423] = 255;
assign img[ 6424] = 221;
assign img[ 6425] = 255;
assign img[ 6426] = 221;
assign img[ 6427] = 255;
assign img[ 6428] = 255;
assign img[ 6429] = 255;
assign img[ 6430] = 239;
assign img[ 6431] = 174;
assign img[ 6432] = 138;
assign img[ 6433] = 238;
assign img[ 6434] = 238;
assign img[ 6435] = 255;
assign img[ 6436] = 255;
assign img[ 6437] = 255;
assign img[ 6438] = 255;
assign img[ 6439] = 239;
assign img[ 6440] = 238;
assign img[ 6441] = 238;
assign img[ 6442] = 238;
assign img[ 6443] = 238;
assign img[ 6444] = 255;
assign img[ 6445] = 254;
assign img[ 6446] = 254;
assign img[ 6447] = 255;
assign img[ 6448] = 255;
assign img[ 6449] = 255;
assign img[ 6450] = 239;
assign img[ 6451] = 238;
assign img[ 6452] = 238;
assign img[ 6453] = 255;
assign img[ 6454] = 255;
assign img[ 6455] = 239;
assign img[ 6456] = 238;
assign img[ 6457] = 238;
assign img[ 6458] = 254;
assign img[ 6459] = 255;
assign img[ 6460] = 255;
assign img[ 6461] = 255;
assign img[ 6462] = 255;
assign img[ 6463] = 255;
assign img[ 6464] = 255;
assign img[ 6465] = 255;
assign img[ 6466] = 255;
assign img[ 6467] = 255;
assign img[ 6468] = 255;
assign img[ 6469] = 255;
assign img[ 6470] = 255;
assign img[ 6471] = 255;
assign img[ 6472] = 255;
assign img[ 6473] = 255;
assign img[ 6474] = 255;
assign img[ 6475] = 255;
assign img[ 6476] = 255;
assign img[ 6477] = 255;
assign img[ 6478] = 238;
assign img[ 6479] = 255;
assign img[ 6480] = 255;
assign img[ 6481] = 255;
assign img[ 6482] = 255;
assign img[ 6483] = 239;
assign img[ 6484] = 238;
assign img[ 6485] = 239;
assign img[ 6486] = 238;
assign img[ 6487] = 238;
assign img[ 6488] = 238;
assign img[ 6489] = 238;
assign img[ 6490] = 238;
assign img[ 6491] = 255;
assign img[ 6492] = 255;
assign img[ 6493] = 255;
assign img[ 6494] = 255;
assign img[ 6495] = 223;
assign img[ 6496] = 204;
assign img[ 6497] = 204;
assign img[ 6498] = 252;
assign img[ 6499] = 255;
assign img[ 6500] = 255;
assign img[ 6501] = 239;
assign img[ 6502] = 254;
assign img[ 6503] = 255;
assign img[ 6504] = 239;
assign img[ 6505] = 238;
assign img[ 6506] = 238;
assign img[ 6507] = 255;
assign img[ 6508] = 239;
assign img[ 6509] = 238;
assign img[ 6510] = 238;
assign img[ 6511] = 238;
assign img[ 6512] = 206;
assign img[ 6513] = 238;
assign img[ 6514] = 238;
assign img[ 6515] = 238;
assign img[ 6516] = 206;
assign img[ 6517] = 238;
assign img[ 6518] = 238;
assign img[ 6519] = 238;
assign img[ 6520] = 238;
assign img[ 6521] = 238;
assign img[ 6522] = 254;
assign img[ 6523] = 255;
assign img[ 6524] = 206;
assign img[ 6525] = 238;
assign img[ 6526] = 238;
assign img[ 6527] = 238;
assign img[ 6528] = 64;
assign img[ 6529] = 68;
assign img[ 6530] = 116;
assign img[ 6531] = 255;
assign img[ 6532] = 238;
assign img[ 6533] = 238;
assign img[ 6534] = 222;
assign img[ 6535] = 255;
assign img[ 6536] = 255;
assign img[ 6537] = 239;
assign img[ 6538] = 238;
assign img[ 6539] = 255;
assign img[ 6540] = 255;
assign img[ 6541] = 255;
assign img[ 6542] = 255;
assign img[ 6543] = 255;
assign img[ 6544] = 239;
assign img[ 6545] = 238;
assign img[ 6546] = 238;
assign img[ 6547] = 255;
assign img[ 6548] = 255;
assign img[ 6549] = 255;
assign img[ 6550] = 239;
assign img[ 6551] = 254;
assign img[ 6552] = 255;
assign img[ 6553] = 207;
assign img[ 6554] = 220;
assign img[ 6555] = 253;
assign img[ 6556] = 255;
assign img[ 6557] = 255;
assign img[ 6558] = 223;
assign img[ 6559] = 205;
assign img[ 6560] = 236;
assign img[ 6561] = 255;
assign img[ 6562] = 255;
assign img[ 6563] = 255;
assign img[ 6564] = 255;
assign img[ 6565] = 255;
assign img[ 6566] = 255;
assign img[ 6567] = 255;
assign img[ 6568] = 238;
assign img[ 6569] = 255;
assign img[ 6570] = 254;
assign img[ 6571] = 255;
assign img[ 6572] = 255;
assign img[ 6573] = 255;
assign img[ 6574] = 255;
assign img[ 6575] = 223;
assign img[ 6576] = 255;
assign img[ 6577] = 239;
assign img[ 6578] = 238;
assign img[ 6579] = 238;
assign img[ 6580] = 206;
assign img[ 6581] = 238;
assign img[ 6582] = 238;
assign img[ 6583] = 254;
assign img[ 6584] = 254;
assign img[ 6585] = 255;
assign img[ 6586] = 222;
assign img[ 6587] = 255;
assign img[ 6588] = 255;
assign img[ 6589] = 255;
assign img[ 6590] = 239;
assign img[ 6591] = 238;
assign img[ 6592] = 238;
assign img[ 6593] = 207;
assign img[ 6594] = 238;
assign img[ 6595] = 238;
assign img[ 6596] = 254;
assign img[ 6597] = 255;
assign img[ 6598] = 255;
assign img[ 6599] = 255;
assign img[ 6600] = 255;
assign img[ 6601] = 255;
assign img[ 6602] = 255;
assign img[ 6603] = 223;
assign img[ 6604] = 221;
assign img[ 6605] = 255;
assign img[ 6606] = 255;
assign img[ 6607] = 255;
assign img[ 6608] = 207;
assign img[ 6609] = 238;
assign img[ 6610] = 238;
assign img[ 6611] = 238;
assign img[ 6612] = 238;
assign img[ 6613] = 255;
assign img[ 6614] = 255;
assign img[ 6615] = 255;
assign img[ 6616] = 255;
assign img[ 6617] = 255;
assign img[ 6618] = 255;
assign img[ 6619] = 255;
assign img[ 6620] = 255;
assign img[ 6621] = 255;
assign img[ 6622] = 255;
assign img[ 6623] = 255;
assign img[ 6624] = 155;
assign img[ 6625] = 223;
assign img[ 6626] = 255;
assign img[ 6627] = 255;
assign img[ 6628] = 255;
assign img[ 6629] = 223;
assign img[ 6630] = 221;
assign img[ 6631] = 253;
assign img[ 6632] = 255;
assign img[ 6633] = 255;
assign img[ 6634] = 255;
assign img[ 6635] = 255;
assign img[ 6636] = 255;
assign img[ 6637] = 255;
assign img[ 6638] = 255;
assign img[ 6639] = 255;
assign img[ 6640] = 221;
assign img[ 6641] = 255;
assign img[ 6642] = 255;
assign img[ 6643] = 255;
assign img[ 6644] = 255;
assign img[ 6645] = 255;
assign img[ 6646] = 255;
assign img[ 6647] = 255;
assign img[ 6648] = 255;
assign img[ 6649] = 255;
assign img[ 6650] = 255;
assign img[ 6651] = 255;
assign img[ 6652] = 239;
assign img[ 6653] = 255;
assign img[ 6654] = 223;
assign img[ 6655] = 221;
assign img[ 6656] = 96;
assign img[ 6657] = 238;
assign img[ 6658] = 238;
assign img[ 6659] = 238;
assign img[ 6660] = 206;
assign img[ 6661] = 238;
assign img[ 6662] = 206;
assign img[ 6663] = 254;
assign img[ 6664] = 238;
assign img[ 6665] = 255;
assign img[ 6666] = 255;
assign img[ 6667] = 255;
assign img[ 6668] = 204;
assign img[ 6669] = 238;
assign img[ 6670] = 238;
assign img[ 6671] = 238;
assign img[ 6672] = 238;
assign img[ 6673] = 238;
assign img[ 6674] = 238;
assign img[ 6675] = 238;
assign img[ 6676] = 220;
assign img[ 6677] = 221;
assign img[ 6678] = 239;
assign img[ 6679] = 238;
assign img[ 6680] = 238;
assign img[ 6681] = 255;
assign img[ 6682] = 255;
assign img[ 6683] = 255;
assign img[ 6684] = 255;
assign img[ 6685] = 255;
assign img[ 6686] = 255;
assign img[ 6687] = 255;
assign img[ 6688] = 255;
assign img[ 6689] = 255;
assign img[ 6690] = 239;
assign img[ 6691] = 238;
assign img[ 6692] = 238;
assign img[ 6693] = 238;
assign img[ 6694] = 238;
assign img[ 6695] = 238;
assign img[ 6696] = 238;
assign img[ 6697] = 238;
assign img[ 6698] = 255;
assign img[ 6699] = 255;
assign img[ 6700] = 255;
assign img[ 6701] = 223;
assign img[ 6702] = 253;
assign img[ 6703] = 239;
assign img[ 6704] = 254;
assign img[ 6705] = 255;
assign img[ 6706] = 255;
assign img[ 6707] = 255;
assign img[ 6708] = 255;
assign img[ 6709] = 255;
assign img[ 6710] = 255;
assign img[ 6711] = 255;
assign img[ 6712] = 255;
assign img[ 6713] = 255;
assign img[ 6714] = 255;
assign img[ 6715] = 255;
assign img[ 6716] = 255;
assign img[ 6717] = 255;
assign img[ 6718] = 255;
assign img[ 6719] = 255;
assign img[ 6720] = 255;
assign img[ 6721] = 255;
assign img[ 6722] = 255;
assign img[ 6723] = 255;
assign img[ 6724] = 255;
assign img[ 6725] = 255;
assign img[ 6726] = 255;
assign img[ 6727] = 255;
assign img[ 6728] = 255;
assign img[ 6729] = 255;
assign img[ 6730] = 255;
assign img[ 6731] = 255;
assign img[ 6732] = 255;
assign img[ 6733] = 255;
assign img[ 6734] = 254;
assign img[ 6735] = 255;
assign img[ 6736] = 255;
assign img[ 6737] = 255;
assign img[ 6738] = 255;
assign img[ 6739] = 255;
assign img[ 6740] = 238;
assign img[ 6741] = 238;
assign img[ 6742] = 238;
assign img[ 6743] = 254;
assign img[ 6744] = 255;
assign img[ 6745] = 255;
assign img[ 6746] = 255;
assign img[ 6747] = 255;
assign img[ 6748] = 238;
assign img[ 6749] = 255;
assign img[ 6750] = 238;
assign img[ 6751] = 223;
assign img[ 6752] = 221;
assign img[ 6753] = 253;
assign img[ 6754] = 255;
assign img[ 6755] = 255;
assign img[ 6756] = 255;
assign img[ 6757] = 255;
assign img[ 6758] = 187;
assign img[ 6759] = 251;
assign img[ 6760] = 255;
assign img[ 6761] = 255;
assign img[ 6762] = 204;
assign img[ 6763] = 238;
assign img[ 6764] = 222;
assign img[ 6765] = 255;
assign img[ 6766] = 255;
assign img[ 6767] = 255;
assign img[ 6768] = 239;
assign img[ 6769] = 238;
assign img[ 6770] = 238;
assign img[ 6771] = 254;
assign img[ 6772] = 223;
assign img[ 6773] = 205;
assign img[ 6774] = 236;
assign img[ 6775] = 255;
assign img[ 6776] = 255;
assign img[ 6777] = 255;
assign img[ 6778] = 255;
assign img[ 6779] = 207;
assign img[ 6780] = 220;
assign img[ 6781] = 255;
assign img[ 6782] = 255;
assign img[ 6783] = 255;
assign img[ 6784] = 96;
assign img[ 6785] = 207;
assign img[ 6786] = 253;
assign img[ 6787] = 255;
assign img[ 6788] = 239;
assign img[ 6789] = 238;
assign img[ 6790] = 238;
assign img[ 6791] = 238;
assign img[ 6792] = 238;
assign img[ 6793] = 238;
assign img[ 6794] = 238;
assign img[ 6795] = 254;
assign img[ 6796] = 255;
assign img[ 6797] = 255;
assign img[ 6798] = 255;
assign img[ 6799] = 223;
assign img[ 6800] = 253;
assign img[ 6801] = 255;
assign img[ 6802] = 255;
assign img[ 6803] = 255;
assign img[ 6804] = 255;
assign img[ 6805] = 238;
assign img[ 6806] = 238;
assign img[ 6807] = 255;
assign img[ 6808] = 255;
assign img[ 6809] = 255;
assign img[ 6810] = 255;
assign img[ 6811] = 255;
assign img[ 6812] = 255;
assign img[ 6813] = 255;
assign img[ 6814] = 255;
assign img[ 6815] = 255;
assign img[ 6816] = 255;
assign img[ 6817] = 255;
assign img[ 6818] = 255;
assign img[ 6819] = 255;
assign img[ 6820] = 255;
assign img[ 6821] = 255;
assign img[ 6822] = 255;
assign img[ 6823] = 223;
assign img[ 6824] = 239;
assign img[ 6825] = 238;
assign img[ 6826] = 238;
assign img[ 6827] = 238;
assign img[ 6828] = 238;
assign img[ 6829] = 206;
assign img[ 6830] = 252;
assign img[ 6831] = 255;
assign img[ 6832] = 255;
assign img[ 6833] = 255;
assign img[ 6834] = 239;
assign img[ 6835] = 238;
assign img[ 6836] = 238;
assign img[ 6837] = 255;
assign img[ 6838] = 239;
assign img[ 6839] = 238;
assign img[ 6840] = 238;
assign img[ 6841] = 238;
assign img[ 6842] = 254;
assign img[ 6843] = 255;
assign img[ 6844] = 255;
assign img[ 6845] = 255;
assign img[ 6846] = 238;
assign img[ 6847] = 255;
assign img[ 6848] = 255;
assign img[ 6849] = 255;
assign img[ 6850] = 239;
assign img[ 6851] = 255;
assign img[ 6852] = 255;
assign img[ 6853] = 255;
assign img[ 6854] = 255;
assign img[ 6855] = 239;
assign img[ 6856] = 238;
assign img[ 6857] = 239;
assign img[ 6858] = 255;
assign img[ 6859] = 255;
assign img[ 6860] = 255;
assign img[ 6861] = 255;
assign img[ 6862] = 238;
assign img[ 6863] = 255;
assign img[ 6864] = 255;
assign img[ 6865] = 255;
assign img[ 6866] = 255;
assign img[ 6867] = 239;
assign img[ 6868] = 238;
assign img[ 6869] = 238;
assign img[ 6870] = 238;
assign img[ 6871] = 255;
assign img[ 6872] = 255;
assign img[ 6873] = 255;
assign img[ 6874] = 255;
assign img[ 6875] = 255;
assign img[ 6876] = 255;
assign img[ 6877] = 255;
assign img[ 6878] = 255;
assign img[ 6879] = 223;
assign img[ 6880] = 221;
assign img[ 6881] = 253;
assign img[ 6882] = 255;
assign img[ 6883] = 255;
assign img[ 6884] = 255;
assign img[ 6885] = 255;
assign img[ 6886] = 221;
assign img[ 6887] = 255;
assign img[ 6888] = 255;
assign img[ 6889] = 255;
assign img[ 6890] = 255;
assign img[ 6891] = 239;
assign img[ 6892] = 206;
assign img[ 6893] = 238;
assign img[ 6894] = 238;
assign img[ 6895] = 238;
assign img[ 6896] = 254;
assign img[ 6897] = 239;
assign img[ 6898] = 238;
assign img[ 6899] = 238;
assign img[ 6900] = 254;
assign img[ 6901] = 255;
assign img[ 6902] = 255;
assign img[ 6903] = 255;
assign img[ 6904] = 255;
assign img[ 6905] = 255;
assign img[ 6906] = 255;
assign img[ 6907] = 255;
assign img[ 6908] = 238;
assign img[ 6909] = 255;
assign img[ 6910] = 207;
assign img[ 6911] = 238;
assign img[ 6912] = 96;
assign img[ 6913] = 255;
assign img[ 6914] = 255;
assign img[ 6915] = 239;
assign img[ 6916] = 238;
assign img[ 6917] = 238;
assign img[ 6918] = 238;
assign img[ 6919] = 238;
assign img[ 6920] = 238;
assign img[ 6921] = 238;
assign img[ 6922] = 238;
assign img[ 6923] = 254;
assign img[ 6924] = 239;
assign img[ 6925] = 254;
assign img[ 6926] = 221;
assign img[ 6927] = 253;
assign img[ 6928] = 223;
assign img[ 6929] = 221;
assign img[ 6930] = 253;
assign img[ 6931] = 255;
assign img[ 6932] = 255;
assign img[ 6933] = 255;
assign img[ 6934] = 255;
assign img[ 6935] = 255;
assign img[ 6936] = 255;
assign img[ 6937] = 255;
assign img[ 6938] = 221;
assign img[ 6939] = 221;
assign img[ 6940] = 253;
assign img[ 6941] = 255;
assign img[ 6942] = 255;
assign img[ 6943] = 239;
assign img[ 6944] = 220;
assign img[ 6945] = 255;
assign img[ 6946] = 255;
assign img[ 6947] = 255;
assign img[ 6948] = 255;
assign img[ 6949] = 239;
assign img[ 6950] = 238;
assign img[ 6951] = 238;
assign img[ 6952] = 238;
assign img[ 6953] = 238;
assign img[ 6954] = 238;
assign img[ 6955] = 238;
assign img[ 6956] = 238;
assign img[ 6957] = 238;
assign img[ 6958] = 238;
assign img[ 6959] = 255;
assign img[ 6960] = 255;
assign img[ 6961] = 255;
assign img[ 6962] = 255;
assign img[ 6963] = 255;
assign img[ 6964] = 255;
assign img[ 6965] = 255;
assign img[ 6966] = 255;
assign img[ 6967] = 255;
assign img[ 6968] = 255;
assign img[ 6969] = 255;
assign img[ 6970] = 255;
assign img[ 6971] = 255;
assign img[ 6972] = 255;
assign img[ 6973] = 223;
assign img[ 6974] = 255;
assign img[ 6975] = 255;
assign img[ 6976] = 255;
assign img[ 6977] = 255;
assign img[ 6978] = 223;
assign img[ 6979] = 255;
assign img[ 6980] = 255;
assign img[ 6981] = 255;
assign img[ 6982] = 221;
assign img[ 6983] = 205;
assign img[ 6984] = 238;
assign img[ 6985] = 255;
assign img[ 6986] = 255;
assign img[ 6987] = 255;
assign img[ 6988] = 255;
assign img[ 6989] = 255;
assign img[ 6990] = 255;
assign img[ 6991] = 255;
assign img[ 6992] = 255;
assign img[ 6993] = 255;
assign img[ 6994] = 255;
assign img[ 6995] = 255;
assign img[ 6996] = 255;
assign img[ 6997] = 223;
assign img[ 6998] = 236;
assign img[ 6999] = 238;
assign img[ 7000] = 254;
assign img[ 7001] = 255;
assign img[ 7002] = 255;
assign img[ 7003] = 255;
assign img[ 7004] = 255;
assign img[ 7005] = 255;
assign img[ 7006] = 255;
assign img[ 7007] = 255;
assign img[ 7008] = 155;
assign img[ 7009] = 255;
assign img[ 7010] = 255;
assign img[ 7011] = 255;
assign img[ 7012] = 255;
assign img[ 7013] = 255;
assign img[ 7014] = 221;
assign img[ 7015] = 253;
assign img[ 7016] = 255;
assign img[ 7017] = 255;
assign img[ 7018] = 255;
assign img[ 7019] = 255;
assign img[ 7020] = 187;
assign img[ 7021] = 251;
assign img[ 7022] = 251;
assign img[ 7023] = 255;
assign img[ 7024] = 239;
assign img[ 7025] = 255;
assign img[ 7026] = 255;
assign img[ 7027] = 239;
assign img[ 7028] = 238;
assign img[ 7029] = 238;
assign img[ 7030] = 238;
assign img[ 7031] = 238;
assign img[ 7032] = 254;
assign img[ 7033] = 239;
assign img[ 7034] = 238;
assign img[ 7035] = 238;
assign img[ 7036] = 238;
assign img[ 7037] = 238;
assign img[ 7038] = 238;
assign img[ 7039] = 255;
assign img[ 7040] = 96;
assign img[ 7041] = 255;
assign img[ 7042] = 255;
assign img[ 7043] = 207;
assign img[ 7044] = 204;
assign img[ 7045] = 204;
assign img[ 7046] = 220;
assign img[ 7047] = 255;
assign img[ 7048] = 255;
assign img[ 7049] = 255;
assign img[ 7050] = 255;
assign img[ 7051] = 207;
assign img[ 7052] = 236;
assign img[ 7053] = 238;
assign img[ 7054] = 254;
assign img[ 7055] = 239;
assign img[ 7056] = 222;
assign img[ 7057] = 255;
assign img[ 7058] = 255;
assign img[ 7059] = 255;
assign img[ 7060] = 255;
assign img[ 7061] = 255;
assign img[ 7062] = 223;
assign img[ 7063] = 221;
assign img[ 7064] = 236;
assign img[ 7065] = 255;
assign img[ 7066] = 187;
assign img[ 7067] = 255;
assign img[ 7068] = 255;
assign img[ 7069] = 255;
assign img[ 7070] = 239;
assign img[ 7071] = 206;
assign img[ 7072] = 204;
assign img[ 7073] = 253;
assign img[ 7074] = 255;
assign img[ 7075] = 255;
assign img[ 7076] = 255;
assign img[ 7077] = 255;
assign img[ 7078] = 255;
assign img[ 7079] = 255;
assign img[ 7080] = 238;
assign img[ 7081] = 254;
assign img[ 7082] = 238;
assign img[ 7083] = 238;
assign img[ 7084] = 238;
assign img[ 7085] = 238;
assign img[ 7086] = 238;
assign img[ 7087] = 238;
assign img[ 7088] = 238;
assign img[ 7089] = 255;
assign img[ 7090] = 255;
assign img[ 7091] = 223;
assign img[ 7092] = 221;
assign img[ 7093] = 255;
assign img[ 7094] = 255;
assign img[ 7095] = 255;
assign img[ 7096] = 255;
assign img[ 7097] = 255;
assign img[ 7098] = 238;
assign img[ 7099] = 238;
assign img[ 7100] = 254;
assign img[ 7101] = 255;
assign img[ 7102] = 187;
assign img[ 7103] = 255;
assign img[ 7104] = 255;
assign img[ 7105] = 255;
assign img[ 7106] = 255;
assign img[ 7107] = 255;
assign img[ 7108] = 255;
assign img[ 7109] = 255;
assign img[ 7110] = 239;
assign img[ 7111] = 238;
assign img[ 7112] = 238;
assign img[ 7113] = 238;
assign img[ 7114] = 254;
assign img[ 7115] = 255;
assign img[ 7116] = 223;
assign img[ 7117] = 239;
assign img[ 7118] = 238;
assign img[ 7119] = 238;
assign img[ 7120] = 254;
assign img[ 7121] = 255;
assign img[ 7122] = 223;
assign img[ 7123] = 255;
assign img[ 7124] = 255;
assign img[ 7125] = 255;
assign img[ 7126] = 255;
assign img[ 7127] = 255;
assign img[ 7128] = 255;
assign img[ 7129] = 255;
assign img[ 7130] = 255;
assign img[ 7131] = 255;
assign img[ 7132] = 255;
assign img[ 7133] = 255;
assign img[ 7134] = 255;
assign img[ 7135] = 223;
assign img[ 7136] = 253;
assign img[ 7137] = 255;
assign img[ 7138] = 238;
assign img[ 7139] = 238;
assign img[ 7140] = 238;
assign img[ 7141] = 255;
assign img[ 7142] = 204;
assign img[ 7143] = 238;
assign img[ 7144] = 254;
assign img[ 7145] = 255;
assign img[ 7146] = 255;
assign img[ 7147] = 239;
assign img[ 7148] = 174;
assign img[ 7149] = 238;
assign img[ 7150] = 238;
assign img[ 7151] = 206;
assign img[ 7152] = 236;
assign img[ 7153] = 238;
assign img[ 7154] = 254;
assign img[ 7155] = 239;
assign img[ 7156] = 222;
assign img[ 7157] = 204;
assign img[ 7158] = 236;
assign img[ 7159] = 255;
assign img[ 7160] = 255;
assign img[ 7161] = 255;
assign img[ 7162] = 255;
assign img[ 7163] = 238;
assign img[ 7164] = 238;
assign img[ 7165] = 238;
assign img[ 7166] = 238;
assign img[ 7167] = 238;
assign img[ 7168] = 96;
assign img[ 7169] = 223;
assign img[ 7170] = 253;
assign img[ 7171] = 255;
assign img[ 7172] = 223;
assign img[ 7173] = 255;
assign img[ 7174] = 191;
assign img[ 7175] = 170;
assign img[ 7176] = 234;
assign img[ 7177] = 238;
assign img[ 7178] = 238;
assign img[ 7179] = 255;
assign img[ 7180] = 221;
assign img[ 7181] = 253;
assign img[ 7182] = 255;
assign img[ 7183] = 239;
assign img[ 7184] = 238;
assign img[ 7185] = 238;
assign img[ 7186] = 238;
assign img[ 7187] = 142;
assign img[ 7188] = 136;
assign img[ 7189] = 234;
assign img[ 7190] = 206;
assign img[ 7191] = 236;
assign img[ 7192] = 238;
assign img[ 7193] = 238;
assign img[ 7194] = 238;
assign img[ 7195] = 238;
assign img[ 7196] = 238;
assign img[ 7197] = 238;
assign img[ 7198] = 238;
assign img[ 7199] = 206;
assign img[ 7200] = 220;
assign img[ 7201] = 255;
assign img[ 7202] = 255;
assign img[ 7203] = 255;
assign img[ 7204] = 255;
assign img[ 7205] = 255;
assign img[ 7206] = 238;
assign img[ 7207] = 255;
assign img[ 7208] = 238;
assign img[ 7209] = 238;
assign img[ 7210] = 238;
assign img[ 7211] = 238;
assign img[ 7212] = 238;
assign img[ 7213] = 254;
assign img[ 7214] = 255;
assign img[ 7215] = 255;
assign img[ 7216] = 238;
assign img[ 7217] = 238;
assign img[ 7218] = 238;
assign img[ 7219] = 238;
assign img[ 7220] = 238;
assign img[ 7221] = 255;
assign img[ 7222] = 255;
assign img[ 7223] = 255;
assign img[ 7224] = 255;
assign img[ 7225] = 255;
assign img[ 7226] = 190;
assign img[ 7227] = 255;
assign img[ 7228] = 255;
assign img[ 7229] = 255;
assign img[ 7230] = 255;
assign img[ 7231] = 255;
assign img[ 7232] = 255;
assign img[ 7233] = 255;
assign img[ 7234] = 239;
assign img[ 7235] = 238;
assign img[ 7236] = 254;
assign img[ 7237] = 255;
assign img[ 7238] = 255;
assign img[ 7239] = 239;
assign img[ 7240] = 238;
assign img[ 7241] = 238;
assign img[ 7242] = 254;
assign img[ 7243] = 239;
assign img[ 7244] = 254;
assign img[ 7245] = 255;
assign img[ 7246] = 255;
assign img[ 7247] = 255;
assign img[ 7248] = 239;
assign img[ 7249] = 238;
assign img[ 7250] = 238;
assign img[ 7251] = 239;
assign img[ 7252] = 238;
assign img[ 7253] = 238;
assign img[ 7254] = 238;
assign img[ 7255] = 238;
assign img[ 7256] = 238;
assign img[ 7257] = 238;
assign img[ 7258] = 238;
assign img[ 7259] = 238;
assign img[ 7260] = 238;
assign img[ 7261] = 238;
assign img[ 7262] = 254;
assign img[ 7263] = 255;
assign img[ 7264] = 187;
assign img[ 7265] = 171;
assign img[ 7266] = 238;
assign img[ 7267] = 238;
assign img[ 7268] = 238;
assign img[ 7269] = 255;
assign img[ 7270] = 255;
assign img[ 7271] = 255;
assign img[ 7272] = 255;
assign img[ 7273] = 255;
assign img[ 7274] = 238;
assign img[ 7275] = 191;
assign img[ 7276] = 155;
assign img[ 7277] = 251;
assign img[ 7278] = 255;
assign img[ 7279] = 255;
assign img[ 7280] = 255;
assign img[ 7281] = 239;
assign img[ 7282] = 238;
assign img[ 7283] = 206;
assign img[ 7284] = 204;
assign img[ 7285] = 236;
assign img[ 7286] = 238;
assign img[ 7287] = 254;
assign img[ 7288] = 255;
assign img[ 7289] = 238;
assign img[ 7290] = 238;
assign img[ 7291] = 206;
assign img[ 7292] = 238;
assign img[ 7293] = 255;
assign img[ 7294] = 223;
assign img[ 7295] = 255;
assign img[ 7296] = 96;
assign img[ 7297] = 174;
assign img[ 7298] = 234;
assign img[ 7299] = 238;
assign img[ 7300] = 238;
assign img[ 7301] = 255;
assign img[ 7302] = 239;
assign img[ 7303] = 254;
assign img[ 7304] = 255;
assign img[ 7305] = 255;
assign img[ 7306] = 255;
assign img[ 7307] = 255;
assign img[ 7308] = 221;
assign img[ 7309] = 221;
assign img[ 7310] = 236;
assign img[ 7311] = 223;
assign img[ 7312] = 221;
assign img[ 7313] = 204;
assign img[ 7314] = 236;
assign img[ 7315] = 238;
assign img[ 7316] = 110;
assign img[ 7317] = 238;
assign img[ 7318] = 238;
assign img[ 7319] = 255;
assign img[ 7320] = 255;
assign img[ 7321] = 255;
assign img[ 7322] = 236;
assign img[ 7323] = 238;
assign img[ 7324] = 238;
assign img[ 7325] = 238;
assign img[ 7326] = 254;
assign img[ 7327] = 255;
assign img[ 7328] = 187;
assign img[ 7329] = 251;
assign img[ 7330] = 255;
assign img[ 7331] = 255;
assign img[ 7332] = 254;
assign img[ 7333] = 174;
assign img[ 7334] = 170;
assign img[ 7335] = 170;
assign img[ 7336] = 234;
assign img[ 7337] = 238;
assign img[ 7338] = 221;
assign img[ 7339] = 253;
assign img[ 7340] = 255;
assign img[ 7341] = 255;
assign img[ 7342] = 255;
assign img[ 7343] = 255;
assign img[ 7344] = 255;
assign img[ 7345] = 239;
assign img[ 7346] = 220;
assign img[ 7347] = 255;
assign img[ 7348] = 223;
assign img[ 7349] = 255;
assign img[ 7350] = 255;
assign img[ 7351] = 255;
assign img[ 7352] = 255;
assign img[ 7353] = 255;
assign img[ 7354] = 239;
assign img[ 7355] = 238;
assign img[ 7356] = 238;
assign img[ 7357] = 255;
assign img[ 7358] = 220;
assign img[ 7359] = 253;
assign img[ 7360] = 255;
assign img[ 7361] = 255;
assign img[ 7362] = 205;
assign img[ 7363] = 236;
assign img[ 7364] = 238;
assign img[ 7365] = 255;
assign img[ 7366] = 238;
assign img[ 7367] = 238;
assign img[ 7368] = 238;
assign img[ 7369] = 255;
assign img[ 7370] = 238;
assign img[ 7371] = 255;
assign img[ 7372] = 255;
assign img[ 7373] = 255;
assign img[ 7374] = 223;
assign img[ 7375] = 255;
assign img[ 7376] = 255;
assign img[ 7377] = 255;
assign img[ 7378] = 255;
assign img[ 7379] = 255;
assign img[ 7380] = 255;
assign img[ 7381] = 223;
assign img[ 7382] = 221;
assign img[ 7383] = 253;
assign img[ 7384] = 255;
assign img[ 7385] = 255;
assign img[ 7386] = 255;
assign img[ 7387] = 255;
assign img[ 7388] = 254;
assign img[ 7389] = 255;
assign img[ 7390] = 255;
assign img[ 7391] = 207;
assign img[ 7392] = 236;
assign img[ 7393] = 238;
assign img[ 7394] = 238;
assign img[ 7395] = 238;
assign img[ 7396] = 254;
assign img[ 7397] = 223;
assign img[ 7398] = 137;
assign img[ 7399] = 200;
assign img[ 7400] = 236;
assign img[ 7401] = 255;
assign img[ 7402] = 255;
assign img[ 7403] = 255;
assign img[ 7404] = 255;
assign img[ 7405] = 255;
assign img[ 7406] = 255;
assign img[ 7407] = 239;
assign img[ 7408] = 238;
assign img[ 7409] = 238;
assign img[ 7410] = 238;
assign img[ 7411] = 238;
assign img[ 7412] = 204;
assign img[ 7413] = 204;
assign img[ 7414] = 236;
assign img[ 7415] = 238;
assign img[ 7416] = 238;
assign img[ 7417] = 255;
assign img[ 7418] = 238;
assign img[ 7419] = 238;
assign img[ 7420] = 254;
assign img[ 7421] = 255;
assign img[ 7422] = 255;
assign img[ 7423] = 255;
assign img[ 7424] = 96;
assign img[ 7425] = 206;
assign img[ 7426] = 236;
assign img[ 7427] = 255;
assign img[ 7428] = 187;
assign img[ 7429] = 251;
assign img[ 7430] = 207;
assign img[ 7431] = 238;
assign img[ 7432] = 238;
assign img[ 7433] = 238;
assign img[ 7434] = 238;
assign img[ 7435] = 255;
assign img[ 7436] = 221;
assign img[ 7437] = 221;
assign img[ 7438] = 221;
assign img[ 7439] = 255;
assign img[ 7440] = 185;
assign img[ 7441] = 171;
assign img[ 7442] = 170;
assign img[ 7443] = 138;
assign img[ 7444] = 152;
assign img[ 7445] = 233;
assign img[ 7446] = 254;
assign img[ 7447] = 255;
assign img[ 7448] = 187;
assign img[ 7449] = 251;
assign img[ 7450] = 239;
assign img[ 7451] = 238;
assign img[ 7452] = 254;
assign img[ 7453] = 159;
assign img[ 7454] = 204;
assign img[ 7455] = 204;
assign img[ 7456] = 236;
assign img[ 7457] = 238;
assign img[ 7458] = 238;
assign img[ 7459] = 238;
assign img[ 7460] = 238;
assign img[ 7461] = 206;
assign img[ 7462] = 204;
assign img[ 7463] = 204;
assign img[ 7464] = 236;
assign img[ 7465] = 238;
assign img[ 7466] = 222;
assign img[ 7467] = 221;
assign img[ 7468] = 253;
assign img[ 7469] = 255;
assign img[ 7470] = 238;
assign img[ 7471] = 254;
assign img[ 7472] = 255;
assign img[ 7473] = 255;
assign img[ 7474] = 238;
assign img[ 7475] = 206;
assign img[ 7476] = 204;
assign img[ 7477] = 252;
assign img[ 7478] = 223;
assign img[ 7479] = 253;
assign img[ 7480] = 238;
assign img[ 7481] = 239;
assign img[ 7482] = 255;
assign img[ 7483] = 255;
assign img[ 7484] = 254;
assign img[ 7485] = 238;
assign img[ 7486] = 238;
assign img[ 7487] = 255;
assign img[ 7488] = 255;
assign img[ 7489] = 255;
assign img[ 7490] = 255;
assign img[ 7491] = 255;
assign img[ 7492] = 255;
assign img[ 7493] = 239;
assign img[ 7494] = 238;
assign img[ 7495] = 238;
assign img[ 7496] = 238;
assign img[ 7497] = 254;
assign img[ 7498] = 255;
assign img[ 7499] = 255;
assign img[ 7500] = 255;
assign img[ 7501] = 255;
assign img[ 7502] = 239;
assign img[ 7503] = 255;
assign img[ 7504] = 255;
assign img[ 7505] = 255;
assign img[ 7506] = 255;
assign img[ 7507] = 255;
assign img[ 7508] = 255;
assign img[ 7509] = 223;
assign img[ 7510] = 253;
assign img[ 7511] = 255;
assign img[ 7512] = 239;
assign img[ 7513] = 238;
assign img[ 7514] = 204;
assign img[ 7515] = 221;
assign img[ 7516] = 253;
assign img[ 7517] = 255;
assign img[ 7518] = 255;
assign img[ 7519] = 255;
assign img[ 7520] = 255;
assign img[ 7521] = 255;
assign img[ 7522] = 221;
assign img[ 7523] = 253;
assign img[ 7524] = 155;
assign img[ 7525] = 221;
assign img[ 7526] = 236;
assign img[ 7527] = 174;
assign img[ 7528] = 170;
assign img[ 7529] = 170;
assign img[ 7530] = 234;
assign img[ 7531] = 206;
assign img[ 7532] = 136;
assign img[ 7533] = 136;
assign img[ 7534] = 136;
assign img[ 7535] = 170;
assign img[ 7536] = 170;
assign img[ 7537] = 234;
assign img[ 7538] = 238;
assign img[ 7539] = 238;
assign img[ 7540] = 206;
assign img[ 7541] = 238;
assign img[ 7542] = 238;
assign img[ 7543] = 238;
assign img[ 7544] = 238;
assign img[ 7545] = 255;
assign img[ 7546] = 238;
assign img[ 7547] = 238;
assign img[ 7548] = 238;
assign img[ 7549] = 238;
assign img[ 7550] = 254;
assign img[ 7551] = 255;
assign img[ 7552] = 96;
assign img[ 7553] = 255;
assign img[ 7554] = 255;
assign img[ 7555] = 255;
assign img[ 7556] = 239;
assign img[ 7557] = 238;
assign img[ 7558] = 238;
assign img[ 7559] = 238;
assign img[ 7560] = 238;
assign img[ 7561] = 238;
assign img[ 7562] = 254;
assign img[ 7563] = 255;
assign img[ 7564] = 187;
assign img[ 7565] = 187;
assign img[ 7566] = 251;
assign img[ 7567] = 191;
assign img[ 7568] = 137;
assign img[ 7569] = 170;
assign img[ 7570] = 200;
assign img[ 7571] = 137;
assign img[ 7572] = 136;
assign img[ 7573] = 153;
assign img[ 7574] = 153;
assign img[ 7575] = 185;
assign img[ 7576] = 170;
assign img[ 7577] = 186;
assign img[ 7578] = 59;
assign img[ 7579] = 51;
assign img[ 7580] = 17;
assign img[ 7581] = 129;
assign img[ 7582] = 136;
assign img[ 7583] = 232;
assign img[ 7584] = 136;
assign img[ 7585] = 200;
assign img[ 7586] = 236;
assign img[ 7587] = 238;
assign img[ 7588] = 254;
assign img[ 7589] = 255;
assign img[ 7590] = 255;
assign img[ 7591] = 239;
assign img[ 7592] = 238;
assign img[ 7593] = 238;
assign img[ 7594] = 238;
assign img[ 7595] = 238;
assign img[ 7596] = 238;
assign img[ 7597] = 238;
assign img[ 7598] = 238;
assign img[ 7599] = 238;
assign img[ 7600] = 238;
assign img[ 7601] = 255;
assign img[ 7602] = 254;
assign img[ 7603] = 191;
assign img[ 7604] = 155;
assign img[ 7605] = 251;
assign img[ 7606] = 235;
assign img[ 7607] = 255;
assign img[ 7608] = 255;
assign img[ 7609] = 255;
assign img[ 7610] = 255;
assign img[ 7611] = 255;
assign img[ 7612] = 254;
assign img[ 7613] = 255;
assign img[ 7614] = 254;
assign img[ 7615] = 255;
assign img[ 7616] = 255;
assign img[ 7617] = 255;
assign img[ 7618] = 255;
assign img[ 7619] = 255;
assign img[ 7620] = 255;
assign img[ 7621] = 239;
assign img[ 7622] = 238;
assign img[ 7623] = 238;
assign img[ 7624] = 238;
assign img[ 7625] = 255;
assign img[ 7626] = 255;
assign img[ 7627] = 239;
assign img[ 7628] = 204;
assign img[ 7629] = 238;
assign img[ 7630] = 255;
assign img[ 7631] = 255;
assign img[ 7632] = 255;
assign img[ 7633] = 255;
assign img[ 7634] = 223;
assign img[ 7635] = 255;
assign img[ 7636] = 255;
assign img[ 7637] = 255;
assign img[ 7638] = 238;
assign img[ 7639] = 238;
assign img[ 7640] = 206;
assign img[ 7641] = 254;
assign img[ 7642] = 255;
assign img[ 7643] = 255;
assign img[ 7644] = 238;
assign img[ 7645] = 255;
assign img[ 7646] = 255;
assign img[ 7647] = 255;
assign img[ 7648] = 205;
assign img[ 7649] = 238;
assign img[ 7650] = 170;
assign img[ 7651] = 170;
assign img[ 7652] = 170;
assign img[ 7653] = 170;
assign img[ 7654] = 200;
assign img[ 7655] = 141;
assign img[ 7656] = 168;
assign img[ 7657] = 186;
assign img[ 7658] = 187;
assign img[ 7659] = 187;
assign img[ 7660] = 137;
assign img[ 7661] = 153;
assign img[ 7662] = 153;
assign img[ 7663] = 153;
assign img[ 7664] = 136;
assign img[ 7665] = 221;
assign img[ 7666] = 221;
assign img[ 7667] = 191;
assign img[ 7668] = 187;
assign img[ 7669] = 235;
assign img[ 7670] = 238;
assign img[ 7671] = 238;
assign img[ 7672] = 238;
assign img[ 7673] = 238;
assign img[ 7674] = 238;
assign img[ 7675] = 207;
assign img[ 7676] = 220;
assign img[ 7677] = 255;
assign img[ 7678] = 239;
assign img[ 7679] = 238;
assign img[ 7680] = 96;
assign img[ 7681] = 70;
assign img[ 7682] = 116;
assign img[ 7683] = 223;
assign img[ 7684] = 221;
assign img[ 7685] = 221;
assign img[ 7686] = 191;
assign img[ 7687] = 187;
assign img[ 7688] = 251;
assign img[ 7689] = 239;
assign img[ 7690] = 238;
assign img[ 7691] = 170;
assign img[ 7692] = 136;
assign img[ 7693] = 168;
assign img[ 7694] = 170;
assign img[ 7695] = 138;
assign img[ 7696] = 136;
assign img[ 7697] = 138;
assign img[ 7698] = 186;
assign img[ 7699] = 139;
assign img[ 7700] = 152;
assign img[ 7701] = 187;
assign img[ 7702] = 155;
assign img[ 7703] = 185;
assign img[ 7704] = 155;
assign img[ 7705] = 187;
assign img[ 7706] = 43;
assign img[ 7707] = 6;
assign img[ 7708] = 96;
assign img[ 7709] = 162;
assign img[ 7710] = 34;
assign img[ 7711] = 147;
assign img[ 7712] = 49;
assign img[ 7713] = 235;
assign img[ 7714] = 238;
assign img[ 7715] = 238;
assign img[ 7716] = 254;
assign img[ 7717] = 255;
assign img[ 7718] = 255;
assign img[ 7719] = 255;
assign img[ 7720] = 255;
assign img[ 7721] = 255;
assign img[ 7722] = 255;
assign img[ 7723] = 255;
assign img[ 7724] = 255;
assign img[ 7725] = 255;
assign img[ 7726] = 238;
assign img[ 7727] = 255;
assign img[ 7728] = 255;
assign img[ 7729] = 255;
assign img[ 7730] = 255;
assign img[ 7731] = 255;
assign img[ 7732] = 255;
assign img[ 7733] = 255;
assign img[ 7734] = 239;
assign img[ 7735] = 238;
assign img[ 7736] = 238;
assign img[ 7737] = 238;
assign img[ 7738] = 238;
assign img[ 7739] = 238;
assign img[ 7740] = 254;
assign img[ 7741] = 255;
assign img[ 7742] = 221;
assign img[ 7743] = 255;
assign img[ 7744] = 255;
assign img[ 7745] = 255;
assign img[ 7746] = 223;
assign img[ 7747] = 255;
assign img[ 7748] = 223;
assign img[ 7749] = 221;
assign img[ 7750] = 253;
assign img[ 7751] = 255;
assign img[ 7752] = 255;
assign img[ 7753] = 255;
assign img[ 7754] = 255;
assign img[ 7755] = 255;
assign img[ 7756] = 221;
assign img[ 7757] = 253;
assign img[ 7758] = 255;
assign img[ 7759] = 255;
assign img[ 7760] = 239;
assign img[ 7761] = 238;
assign img[ 7762] = 206;
assign img[ 7763] = 238;
assign img[ 7764] = 254;
assign img[ 7765] = 255;
assign img[ 7766] = 255;
assign img[ 7767] = 255;
assign img[ 7768] = 238;
assign img[ 7769] = 254;
assign img[ 7770] = 174;
assign img[ 7771] = 255;
assign img[ 7772] = 238;
assign img[ 7773] = 255;
assign img[ 7774] = 254;
assign img[ 7775] = 174;
assign img[ 7776] = 138;
assign img[ 7777] = 136;
assign img[ 7778] = 236;
assign img[ 7779] = 190;
assign img[ 7780] = 139;
assign img[ 7781] = 140;
assign img[ 7782] = 184;
assign img[ 7783] = 159;
assign img[ 7784] = 153;
assign img[ 7785] = 153;
assign img[ 7786] = 187;
assign img[ 7787] = 251;
assign img[ 7788] = 255;
assign img[ 7789] = 255;
assign img[ 7790] = 187;
assign img[ 7791] = 155;
assign img[ 7792] = 136;
assign img[ 7793] = 136;
assign img[ 7794] = 186;
assign img[ 7795] = 187;
assign img[ 7796] = 153;
assign img[ 7797] = 153;
assign img[ 7798] = 153;
assign img[ 7799] = 255;
assign img[ 7800] = 255;
assign img[ 7801] = 191;
assign img[ 7802] = 187;
assign img[ 7803] = 255;
assign img[ 7804] = 221;
assign img[ 7805] = 253;
assign img[ 7806] = 223;
assign img[ 7807] = 253;
assign img[ 7808] = 80;
assign img[ 7809] = 197;
assign img[ 7810] = 204;
assign img[ 7811] = 238;
assign img[ 7812] = 238;
assign img[ 7813] = 238;
assign img[ 7814] = 206;
assign img[ 7815] = 204;
assign img[ 7816] = 236;
assign img[ 7817] = 255;
assign img[ 7818] = 255;
assign img[ 7819] = 137;
assign img[ 7820] = 153;
assign img[ 7821] = 153;
assign img[ 7822] = 153;
assign img[ 7823] = 137;
assign img[ 7824] = 248;
assign img[ 7825] = 191;
assign img[ 7826] = 171;
assign img[ 7827] = 138;
assign img[ 7828] = 136;
assign img[ 7829] = 185;
assign img[ 7830] = 155;
assign img[ 7831] = 185;
assign img[ 7832] = 170;
assign img[ 7833] = 186;
assign img[ 7834] = 42;
assign img[ 7835] = 66;
assign img[ 7836] = 184;
assign img[ 7837] = 155;
assign img[ 7838] = 136;
assign img[ 7839] = 136;
assign img[ 7840] = 24;
assign img[ 7841] = 177;
assign img[ 7842] = 234;
assign img[ 7843] = 238;
assign img[ 7844] = 238;
assign img[ 7845] = 158;
assign img[ 7846] = 249;
assign img[ 7847] = 221;
assign img[ 7848] = 253;
assign img[ 7849] = 255;
assign img[ 7850] = 239;
assign img[ 7851] = 238;
assign img[ 7852] = 238;
assign img[ 7853] = 238;
assign img[ 7854] = 238;
assign img[ 7855] = 255;
assign img[ 7856] = 255;
assign img[ 7857] = 255;
assign img[ 7858] = 239;
assign img[ 7859] = 238;
assign img[ 7860] = 220;
assign img[ 7861] = 253;
assign img[ 7862] = 255;
assign img[ 7863] = 255;
assign img[ 7864] = 255;
assign img[ 7865] = 223;
assign img[ 7866] = 204;
assign img[ 7867] = 238;
assign img[ 7868] = 238;
assign img[ 7869] = 238;
assign img[ 7870] = 238;
assign img[ 7871] = 238;
assign img[ 7872] = 238;
assign img[ 7873] = 255;
assign img[ 7874] = 255;
assign img[ 7875] = 255;
assign img[ 7876] = 255;
assign img[ 7877] = 238;
assign img[ 7878] = 238;
assign img[ 7879] = 238;
assign img[ 7880] = 238;
assign img[ 7881] = 238;
assign img[ 7882] = 238;
assign img[ 7883] = 223;
assign img[ 7884] = 221;
assign img[ 7885] = 253;
assign img[ 7886] = 191;
assign img[ 7887] = 187;
assign img[ 7888] = 219;
assign img[ 7889] = 255;
assign img[ 7890] = 255;
assign img[ 7891] = 255;
assign img[ 7892] = 255;
assign img[ 7893] = 255;
assign img[ 7894] = 238;
assign img[ 7895] = 238;
assign img[ 7896] = 206;
assign img[ 7897] = 223;
assign img[ 7898] = 204;
assign img[ 7899] = 253;
assign img[ 7900] = 238;
assign img[ 7901] = 239;
assign img[ 7902] = 238;
assign img[ 7903] = 174;
assign img[ 7904] = 234;
assign img[ 7905] = 238;
assign img[ 7906] = 136;
assign img[ 7907] = 168;
assign img[ 7908] = 202;
assign img[ 7909] = 140;
assign img[ 7910] = 200;
assign img[ 7911] = 205;
assign img[ 7912] = 221;
assign img[ 7913] = 221;
assign img[ 7914] = 221;
assign img[ 7915] = 157;
assign img[ 7916] = 251;
assign img[ 7917] = 191;
assign img[ 7918] = 138;
assign img[ 7919] = 153;
assign img[ 7920] = 153;
assign img[ 7921] = 157;
assign img[ 7922] = 153;
assign img[ 7923] = 153;
assign img[ 7924] = 137;
assign img[ 7925] = 136;
assign img[ 7926] = 168;
assign img[ 7927] = 234;
assign img[ 7928] = 222;
assign img[ 7929] = 221;
assign img[ 7930] = 236;
assign img[ 7931] = 222;
assign img[ 7932] = 236;
assign img[ 7933] = 255;
assign img[ 7934] = 255;
assign img[ 7935] = 255;
assign img[ 7936] = 96;
assign img[ 7937] = 206;
assign img[ 7938] = 236;
assign img[ 7939] = 238;
assign img[ 7940] = 206;
assign img[ 7941] = 221;
assign img[ 7942] = 221;
assign img[ 7943] = 253;
assign img[ 7944] = 255;
assign img[ 7945] = 239;
assign img[ 7946] = 222;
assign img[ 7947] = 153;
assign img[ 7948] = 249;
assign img[ 7949] = 191;
assign img[ 7950] = 170;
assign img[ 7951] = 138;
assign img[ 7952] = 136;
assign img[ 7953] = 152;
assign img[ 7954] = 153;
assign img[ 7955] = 153;
assign img[ 7956] = 153;
assign img[ 7957] = 153;
assign img[ 7958] = 153;
assign img[ 7959] = 185;
assign img[ 7960] = 187;
assign img[ 7961] = 187;
assign img[ 7962] = 43;
assign img[ 7963] = 34;
assign img[ 7964] = 16;
assign img[ 7965] = 179;
assign img[ 7966] = 138;
assign img[ 7967] = 235;
assign img[ 7968] = 255;
assign img[ 7969] = 255;
assign img[ 7970] = 255;
assign img[ 7971] = 255;
assign img[ 7972] = 255;
assign img[ 7973] = 255;
assign img[ 7974] = 255;
assign img[ 7975] = 255;
assign img[ 7976] = 255;
assign img[ 7977] = 255;
assign img[ 7978] = 239;
assign img[ 7979] = 255;
assign img[ 7980] = 255;
assign img[ 7981] = 255;
assign img[ 7982] = 255;
assign img[ 7983] = 239;
assign img[ 7984] = 238;
assign img[ 7985] = 238;
assign img[ 7986] = 220;
assign img[ 7987] = 221;
assign img[ 7988] = 221;
assign img[ 7989] = 205;
assign img[ 7990] = 221;
assign img[ 7991] = 205;
assign img[ 7992] = 204;
assign img[ 7993] = 236;
assign img[ 7994] = 238;
assign img[ 7995] = 206;
assign img[ 7996] = 204;
assign img[ 7997] = 204;
assign img[ 7998] = 236;
assign img[ 7999] = 255;
assign img[ 8000] = 255;
assign img[ 8001] = 255;
assign img[ 8002] = 255;
assign img[ 8003] = 239;
assign img[ 8004] = 206;
assign img[ 8005] = 221;
assign img[ 8006] = 253;
assign img[ 8007] = 223;
assign img[ 8008] = 236;
assign img[ 8009] = 238;
assign img[ 8010] = 238;
assign img[ 8011] = 238;
assign img[ 8012] = 220;
assign img[ 8013] = 253;
assign img[ 8014] = 255;
assign img[ 8015] = 255;
assign img[ 8016] = 255;
assign img[ 8017] = 255;
assign img[ 8018] = 255;
assign img[ 8019] = 255;
assign img[ 8020] = 255;
assign img[ 8021] = 255;
assign img[ 8022] = 238;
assign img[ 8023] = 238;
assign img[ 8024] = 238;
assign img[ 8025] = 255;
assign img[ 8026] = 254;
assign img[ 8027] = 238;
assign img[ 8028] = 238;
assign img[ 8029] = 238;
assign img[ 8030] = 254;
assign img[ 8031] = 255;
assign img[ 8032] = 239;
assign img[ 8033] = 238;
assign img[ 8034] = 170;
assign img[ 8035] = 170;
assign img[ 8036] = 138;
assign img[ 8037] = 136;
assign img[ 8038] = 168;
assign img[ 8039] = 187;
assign img[ 8040] = 187;
assign img[ 8041] = 155;
assign img[ 8042] = 153;
assign img[ 8043] = 155;
assign img[ 8044] = 137;
assign img[ 8045] = 136;
assign img[ 8046] = 136;
assign img[ 8047] = 153;
assign img[ 8048] = 152;
assign img[ 8049] = 153;
assign img[ 8050] = 169;
assign img[ 8051] = 170;
assign img[ 8052] = 170;
assign img[ 8053] = 170;
assign img[ 8054] = 170;
assign img[ 8055] = 234;
assign img[ 8056] = 238;
assign img[ 8057] = 239;
assign img[ 8058] = 238;
assign img[ 8059] = 255;
assign img[ 8060] = 255;
assign img[ 8061] = 255;
assign img[ 8062] = 255;
assign img[ 8063] = 255;
assign img[ 8064] = 0;
assign img[ 8065] = 136;
assign img[ 8066] = 168;
assign img[ 8067] = 170;
assign img[ 8068] = 186;
assign img[ 8069] = 171;
assign img[ 8070] = 251;
assign img[ 8071] = 255;
assign img[ 8072] = 223;
assign img[ 8073] = 221;
assign img[ 8074] = 221;
assign img[ 8075] = 157;
assign img[ 8076] = 153;
assign img[ 8077] = 153;
assign img[ 8078] = 136;
assign img[ 8079] = 136;
assign img[ 8080] = 136;
assign img[ 8081] = 136;
assign img[ 8082] = 168;
assign img[ 8083] = 138;
assign img[ 8084] = 136;
assign img[ 8085] = 185;
assign img[ 8086] = 155;
assign img[ 8087] = 185;
assign img[ 8088] = 138;
assign img[ 8089] = 136;
assign img[ 8090] = 24;
assign img[ 8091] = 17;
assign img[ 8092] = 32;
assign img[ 8093] = 170;
assign img[ 8094] = 138;
assign img[ 8095] = 168;
assign img[ 8096] = 186;
assign img[ 8097] = 239;
assign img[ 8098] = 238;
assign img[ 8099] = 238;
assign img[ 8100] = 174;
assign img[ 8101] = 254;
assign img[ 8102] = 255;
assign img[ 8103] = 254;
assign img[ 8104] = 238;
assign img[ 8105] = 255;
assign img[ 8106] = 255;
assign img[ 8107] = 255;
assign img[ 8108] = 254;
assign img[ 8109] = 255;
assign img[ 8110] = 254;
assign img[ 8111] = 255;
assign img[ 8112] = 255;
assign img[ 8113] = 239;
assign img[ 8114] = 238;
assign img[ 8115] = 222;
assign img[ 8116] = 157;
assign img[ 8117] = 255;
assign img[ 8118] = 255;
assign img[ 8119] = 255;
assign img[ 8120] = 191;
assign img[ 8121] = 187;
assign img[ 8122] = 187;
assign img[ 8123] = 251;
assign img[ 8124] = 255;
assign img[ 8125] = 255;
assign img[ 8126] = 255;
assign img[ 8127] = 255;
assign img[ 8128] = 255;
assign img[ 8129] = 255;
assign img[ 8130] = 255;
assign img[ 8131] = 255;
assign img[ 8132] = 255;
assign img[ 8133] = 191;
assign img[ 8134] = 187;
assign img[ 8135] = 187;
assign img[ 8136] = 251;
assign img[ 8137] = 255;
assign img[ 8138] = 255;
assign img[ 8139] = 187;
assign img[ 8140] = 187;
assign img[ 8141] = 255;
assign img[ 8142] = 191;
assign img[ 8143] = 255;
assign img[ 8144] = 223;
assign img[ 8145] = 255;
assign img[ 8146] = 191;
assign img[ 8147] = 255;
assign img[ 8148] = 255;
assign img[ 8149] = 239;
assign img[ 8150] = 238;
assign img[ 8151] = 238;
assign img[ 8152] = 254;
assign img[ 8153] = 255;
assign img[ 8154] = 255;
assign img[ 8155] = 255;
assign img[ 8156] = 255;
assign img[ 8157] = 255;
assign img[ 8158] = 223;
assign img[ 8159] = 255;
assign img[ 8160] = 255;
assign img[ 8161] = 239;
assign img[ 8162] = 254;
assign img[ 8163] = 255;
assign img[ 8164] = 139;
assign img[ 8165] = 136;
assign img[ 8166] = 168;
assign img[ 8167] = 155;
assign img[ 8168] = 249;
assign img[ 8169] = 255;
assign img[ 8170] = 153;
assign img[ 8171] = 153;
assign img[ 8172] = 249;
assign img[ 8173] = 255;
assign img[ 8174] = 155;
assign img[ 8175] = 153;
assign img[ 8176] = 136;
assign img[ 8177] = 152;
assign img[ 8178] = 251;
assign img[ 8179] = 239;
assign img[ 8180] = 170;
assign img[ 8181] = 186;
assign img[ 8182] = 187;
assign img[ 8183] = 155;
assign img[ 8184] = 249;
assign img[ 8185] = 255;
assign img[ 8186] = 137;
assign img[ 8187] = 136;
assign img[ 8188] = 249;
assign img[ 8189] = 255;
assign img[ 8190] = 191;
assign img[ 8191] = 255;
assign img[ 8192] = 16;
assign img[ 8193] = 185;
assign img[ 8194] = 251;
assign img[ 8195] = 223;
assign img[ 8196] = 205;
assign img[ 8197] = 204;
assign img[ 8198] = 220;
assign img[ 8199] = 221;
assign img[ 8200] = 221;
assign img[ 8201] = 223;
assign img[ 8202] = 221;
assign img[ 8203] = 205;
assign img[ 8204] = 152;
assign img[ 8205] = 153;
assign img[ 8206] = 153;
assign img[ 8207] = 153;
assign img[ 8208] = 153;
assign img[ 8209] = 153;
assign img[ 8210] = 153;
assign img[ 8211] = 136;
assign img[ 8212] = 136;
assign img[ 8213] = 168;
assign img[ 8214] = 154;
assign img[ 8215] = 153;
assign img[ 8216] = 136;
assign img[ 8217] = 168;
assign img[ 8218] = 42;
assign img[ 8219] = 34;
assign img[ 8220] = 144;
assign img[ 8221] = 153;
assign img[ 8222] = 153;
assign img[ 8223] = 185;
assign img[ 8224] = 187;
assign img[ 8225] = 223;
assign img[ 8226] = 236;
assign img[ 8227] = 238;
assign img[ 8228] = 238;
assign img[ 8229] = 238;
assign img[ 8230] = 238;
assign img[ 8231] = 238;
assign img[ 8232] = 238;
assign img[ 8233] = 238;
assign img[ 8234] = 238;
assign img[ 8235] = 238;
assign img[ 8236] = 254;
assign img[ 8237] = 239;
assign img[ 8238] = 254;
assign img[ 8239] = 255;
assign img[ 8240] = 171;
assign img[ 8241] = 206;
assign img[ 8242] = 204;
assign img[ 8243] = 157;
assign img[ 8244] = 169;
assign img[ 8245] = 234;
assign img[ 8246] = 238;
assign img[ 8247] = 238;
assign img[ 8248] = 254;
assign img[ 8249] = 255;
assign img[ 8250] = 255;
assign img[ 8251] = 255;
assign img[ 8252] = 255;
assign img[ 8253] = 255;
assign img[ 8254] = 255;
assign img[ 8255] = 255;
assign img[ 8256] = 255;
assign img[ 8257] = 255;
assign img[ 8258] = 223;
assign img[ 8259] = 221;
assign img[ 8260] = 253;
assign img[ 8261] = 207;
assign img[ 8262] = 236;
assign img[ 8263] = 238;
assign img[ 8264] = 254;
assign img[ 8265] = 255;
assign img[ 8266] = 255;
assign img[ 8267] = 191;
assign img[ 8268] = 170;
assign img[ 8269] = 170;
assign img[ 8270] = 234;
assign img[ 8271] = 238;
assign img[ 8272] = 222;
assign img[ 8273] = 255;
assign img[ 8274] = 187;
assign img[ 8275] = 187;
assign img[ 8276] = 251;
assign img[ 8277] = 255;
assign img[ 8278] = 255;
assign img[ 8279] = 255;
assign img[ 8280] = 255;
assign img[ 8281] = 255;
assign img[ 8282] = 255;
assign img[ 8283] = 255;
assign img[ 8284] = 255;
assign img[ 8285] = 255;
assign img[ 8286] = 207;
assign img[ 8287] = 204;
assign img[ 8288] = 236;
assign img[ 8289] = 142;
assign img[ 8290] = 232;
assign img[ 8291] = 170;
assign img[ 8292] = 170;
assign img[ 8293] = 138;
assign img[ 8294] = 184;
assign img[ 8295] = 191;
assign img[ 8296] = 201;
assign img[ 8297] = 138;
assign img[ 8298] = 186;
assign img[ 8299] = 155;
assign img[ 8300] = 153;
assign img[ 8301] = 169;
assign img[ 8302] = 152;
assign img[ 8303] = 137;
assign img[ 8304] = 136;
assign img[ 8305] = 136;
assign img[ 8306] = 136;
assign img[ 8307] = 136;
assign img[ 8308] = 136;
assign img[ 8309] = 153;
assign img[ 8310] = 153;
assign img[ 8311] = 185;
assign img[ 8312] = 187;
assign img[ 8313] = 191;
assign img[ 8314] = 187;
assign img[ 8315] = 137;
assign img[ 8316] = 200;
assign img[ 8317] = 253;
assign img[ 8318] = 175;
assign img[ 8319] = 170;
assign img[ 8320] = 64;
assign img[ 8321] = 68;
assign img[ 8322] = 100;
assign img[ 8323] = 255;
assign img[ 8324] = 255;
assign img[ 8325] = 205;
assign img[ 8326] = 204;
assign img[ 8327] = 221;
assign img[ 8328] = 221;
assign img[ 8329] = 205;
assign img[ 8330] = 220;
assign img[ 8331] = 205;
assign img[ 8332] = 136;
assign img[ 8333] = 153;
assign img[ 8334] = 153;
assign img[ 8335] = 153;
assign img[ 8336] = 136;
assign img[ 8337] = 152;
assign img[ 8338] = 137;
assign img[ 8339] = 136;
assign img[ 8340] = 152;
assign img[ 8341] = 153;
assign img[ 8342] = 153;
assign img[ 8343] = 153;
assign img[ 8344] = 153;
assign img[ 8345] = 185;
assign img[ 8346] = 27;
assign img[ 8347] = 17;
assign img[ 8348] = 17;
assign img[ 8349] = 153;
assign img[ 8350] = 153;
assign img[ 8351] = 185;
assign img[ 8352] = 187;
assign img[ 8353] = 187;
assign img[ 8354] = 187;
assign img[ 8355] = 255;
assign img[ 8356] = 239;
assign img[ 8357] = 238;
assign img[ 8358] = 254;
assign img[ 8359] = 255;
assign img[ 8360] = 255;
assign img[ 8361] = 255;
assign img[ 8362] = 255;
assign img[ 8363] = 255;
assign img[ 8364] = 255;
assign img[ 8365] = 191;
assign img[ 8366] = 221;
assign img[ 8367] = 157;
assign img[ 8368] = 249;
assign img[ 8369] = 239;
assign img[ 8370] = 204;
assign img[ 8371] = 220;
assign img[ 8372] = 205;
assign img[ 8373] = 236;
assign img[ 8374] = 238;
assign img[ 8375] = 238;
assign img[ 8376] = 254;
assign img[ 8377] = 255;
assign img[ 8378] = 223;
assign img[ 8379] = 221;
assign img[ 8380] = 221;
assign img[ 8381] = 221;
assign img[ 8382] = 205;
assign img[ 8383] = 140;
assign img[ 8384] = 152;
assign img[ 8385] = 251;
assign img[ 8386] = 255;
assign img[ 8387] = 207;
assign img[ 8388] = 236;
assign img[ 8389] = 238;
assign img[ 8390] = 220;
assign img[ 8391] = 255;
assign img[ 8392] = 255;
assign img[ 8393] = 255;
assign img[ 8394] = 238;
assign img[ 8395] = 255;
assign img[ 8396] = 238;
assign img[ 8397] = 205;
assign img[ 8398] = 221;
assign img[ 8399] = 253;
assign img[ 8400] = 159;
assign img[ 8401] = 221;
assign img[ 8402] = 221;
assign img[ 8403] = 157;
assign img[ 8404] = 217;
assign img[ 8405] = 221;
assign img[ 8406] = 255;
assign img[ 8407] = 255;
assign img[ 8408] = 255;
assign img[ 8409] = 255;
assign img[ 8410] = 221;
assign img[ 8411] = 221;
assign img[ 8412] = 236;
assign img[ 8413] = 254;
assign img[ 8414] = 255;
assign img[ 8415] = 255;
assign img[ 8416] = 255;
assign img[ 8417] = 255;
assign img[ 8418] = 153;
assign img[ 8419] = 153;
assign img[ 8420] = 137;
assign img[ 8421] = 136;
assign img[ 8422] = 184;
assign img[ 8423] = 159;
assign img[ 8424] = 185;
assign img[ 8425] = 187;
assign img[ 8426] = 153;
assign img[ 8427] = 187;
assign img[ 8428] = 153;
assign img[ 8429] = 153;
assign img[ 8430] = 136;
assign img[ 8431] = 136;
assign img[ 8432] = 136;
assign img[ 8433] = 136;
assign img[ 8434] = 168;
assign img[ 8435] = 187;
assign img[ 8436] = 170;
assign img[ 8437] = 136;
assign img[ 8438] = 136;
assign img[ 8439] = 232;
assign img[ 8440] = 206;
assign img[ 8441] = 253;
assign img[ 8442] = 127;
assign img[ 8443] = 223;
assign img[ 8444] = 253;
assign img[ 8445] = 255;
assign img[ 8446] = 223;
assign img[ 8447] = 221;
assign img[ 8448] = 96;
assign img[ 8449] = 223;
assign img[ 8450] = 253;
assign img[ 8451] = 255;
assign img[ 8452] = 187;
assign img[ 8453] = 187;
assign img[ 8454] = 170;
assign img[ 8455] = 187;
assign img[ 8456] = 234;
assign img[ 8457] = 239;
assign img[ 8458] = 221;
assign img[ 8459] = 221;
assign img[ 8460] = 153;
assign img[ 8461] = 153;
assign img[ 8462] = 153;
assign img[ 8463] = 137;
assign img[ 8464] = 136;
assign img[ 8465] = 136;
assign img[ 8466] = 152;
assign img[ 8467] = 139;
assign img[ 8468] = 168;
assign img[ 8469] = 186;
assign img[ 8470] = 187;
assign img[ 8471] = 191;
assign img[ 8472] = 170;
assign img[ 8473] = 187;
assign img[ 8474] = 43;
assign img[ 8475] = 3;
assign img[ 8476] = 224;
assign img[ 8477] = 238;
assign img[ 8478] = 170;
assign img[ 8479] = 170;
assign img[ 8480] = 186;
assign img[ 8481] = 187;
assign img[ 8482] = 251;
assign img[ 8483] = 255;
assign img[ 8484] = 255;
assign img[ 8485] = 255;
assign img[ 8486] = 255;
assign img[ 8487] = 255;
assign img[ 8488] = 238;
assign img[ 8489] = 238;
assign img[ 8490] = 238;
assign img[ 8491] = 238;
assign img[ 8492] = 238;
assign img[ 8493] = 238;
assign img[ 8494] = 204;
assign img[ 8495] = 174;
assign img[ 8496] = 238;
assign img[ 8497] = 238;
assign img[ 8498] = 204;
assign img[ 8499] = 238;
assign img[ 8500] = 238;
assign img[ 8501] = 238;
assign img[ 8502] = 238;
assign img[ 8503] = 238;
assign img[ 8504] = 254;
assign img[ 8505] = 255;
assign img[ 8506] = 223;
assign img[ 8507] = 255;
assign img[ 8508] = 238;
assign img[ 8509] = 222;
assign img[ 8510] = 205;
assign img[ 8511] = 254;
assign img[ 8512] = 239;
assign img[ 8513] = 238;
assign img[ 8514] = 170;
assign img[ 8515] = 238;
assign img[ 8516] = 238;
assign img[ 8517] = 255;
assign img[ 8518] = 255;
assign img[ 8519] = 207;
assign img[ 8520] = 252;
assign img[ 8521] = 255;
assign img[ 8522] = 255;
assign img[ 8523] = 223;
assign img[ 8524] = 253;
assign img[ 8525] = 239;
assign img[ 8526] = 254;
assign img[ 8527] = 239;
assign img[ 8528] = 206;
assign img[ 8529] = 204;
assign img[ 8530] = 220;
assign img[ 8531] = 221;
assign img[ 8532] = 253;
assign img[ 8533] = 255;
assign img[ 8534] = 238;
assign img[ 8535] = 238;
assign img[ 8536] = 238;
assign img[ 8537] = 238;
assign img[ 8538] = 238;
assign img[ 8539] = 238;
assign img[ 8540] = 238;
assign img[ 8541] = 238;
assign img[ 8542] = 255;
assign img[ 8543] = 255;
assign img[ 8544] = 239;
assign img[ 8545] = 174;
assign img[ 8546] = 170;
assign img[ 8547] = 206;
assign img[ 8548] = 204;
assign img[ 8549] = 140;
assign img[ 8550] = 200;
assign img[ 8551] = 157;
assign img[ 8552] = 137;
assign img[ 8553] = 174;
assign img[ 8554] = 170;
assign img[ 8555] = 171;
assign img[ 8556] = 139;
assign img[ 8557] = 170;
assign img[ 8558] = 138;
assign img[ 8559] = 153;
assign img[ 8560] = 153;
assign img[ 8561] = 136;
assign img[ 8562] = 136;
assign img[ 8563] = 153;
assign img[ 8564] = 136;
assign img[ 8565] = 136;
assign img[ 8566] = 200;
assign img[ 8567] = 220;
assign img[ 8568] = 189;
assign img[ 8569] = 187;
assign img[ 8570] = 43;
assign img[ 8571] = 34;
assign img[ 8572] = 178;
assign img[ 8573] = 171;
assign img[ 8574] = 250;
assign img[ 8575] = 255;
assign img[ 8576] = 96;
assign img[ 8577] = 238;
assign img[ 8578] = 254;
assign img[ 8579] = 239;
assign img[ 8580] = 238;
assign img[ 8581] = 142;
assign img[ 8582] = 200;
assign img[ 8583] = 204;
assign img[ 8584] = 168;
assign img[ 8585] = 170;
assign img[ 8586] = 186;
assign img[ 8587] = 171;
assign img[ 8588] = 170;
assign img[ 8589] = 170;
assign img[ 8590] = 187;
assign img[ 8591] = 139;
assign img[ 8592] = 136;
assign img[ 8593] = 152;
assign img[ 8594] = 249;
assign img[ 8595] = 255;
assign img[ 8596] = 191;
assign img[ 8597] = 187;
assign img[ 8598] = 187;
assign img[ 8599] = 171;
assign img[ 8600] = 170;
assign img[ 8601] = 170;
assign img[ 8602] = 42;
assign img[ 8603] = 34;
assign img[ 8604] = 16;
assign img[ 8605] = 145;
assign img[ 8606] = 139;
assign img[ 8607] = 216;
assign img[ 8608] = 51;
assign img[ 8609] = 51;
assign img[ 8610] = 211;
assign img[ 8611] = 255;
assign img[ 8612] = 191;
assign img[ 8613] = 171;
assign img[ 8614] = 234;
assign img[ 8615] = 239;
assign img[ 8616] = 238;
assign img[ 8617] = 238;
assign img[ 8618] = 238;
assign img[ 8619] = 238;
assign img[ 8620] = 238;
assign img[ 8621] = 238;
assign img[ 8622] = 186;
assign img[ 8623] = 255;
assign img[ 8624] = 255;
assign img[ 8625] = 255;
assign img[ 8626] = 223;
assign img[ 8627] = 255;
assign img[ 8628] = 255;
assign img[ 8629] = 255;
assign img[ 8630] = 255;
assign img[ 8631] = 255;
assign img[ 8632] = 239;
assign img[ 8633] = 238;
assign img[ 8634] = 206;
assign img[ 8635] = 238;
assign img[ 8636] = 238;
assign img[ 8637] = 239;
assign img[ 8638] = 204;
assign img[ 8639] = 220;
assign img[ 8640] = 221;
assign img[ 8641] = 221;
assign img[ 8642] = 221;
assign img[ 8643] = 189;
assign img[ 8644] = 251;
assign img[ 8645] = 239;
assign img[ 8646] = 238;
assign img[ 8647] = 239;
assign img[ 8648] = 255;
assign img[ 8649] = 255;
assign img[ 8650] = 187;
assign img[ 8651] = 171;
assign img[ 8652] = 186;
assign img[ 8653] = 159;
assign img[ 8654] = 251;
assign img[ 8655] = 223;
assign img[ 8656] = 137;
assign img[ 8657] = 136;
assign img[ 8658] = 186;
assign img[ 8659] = 187;
assign img[ 8660] = 234;
assign img[ 8661] = 238;
assign img[ 8662] = 238;
assign img[ 8663] = 238;
assign img[ 8664] = 238;
assign img[ 8665] = 238;
assign img[ 8666] = 254;
assign img[ 8667] = 223;
assign img[ 8668] = 253;
assign img[ 8669] = 207;
assign img[ 8670] = 172;
assign img[ 8671] = 238;
assign img[ 8672] = 110;
assign img[ 8673] = 151;
assign img[ 8674] = 17;
assign img[ 8675] = 145;
assign img[ 8676] = 145;
assign img[ 8677] = 253;
assign img[ 8678] = 255;
assign img[ 8679] = 191;
assign img[ 8680] = 170;
assign img[ 8681] = 186;
assign img[ 8682] = 171;
assign img[ 8683] = 186;
assign img[ 8684] = 170;
assign img[ 8685] = 136;
assign img[ 8686] = 136;
assign img[ 8687] = 137;
assign img[ 8688] = 137;
assign img[ 8689] = 136;
assign img[ 8690] = 136;
assign img[ 8691] = 152;
assign img[ 8692] = 153;
assign img[ 8693] = 153;
assign img[ 8694] = 185;
assign img[ 8695] = 170;
assign img[ 8696] = 138;
assign img[ 8697] = 136;
assign img[ 8698] = 152;
assign img[ 8699] = 169;
assign img[ 8700] = 202;
assign img[ 8701] = 204;
assign img[ 8702] = 221;
assign img[ 8703] = 255;
assign img[ 8704] = 96;
assign img[ 8705] = 206;
assign img[ 8706] = 220;
assign img[ 8707] = 207;
assign img[ 8708] = 132;
assign img[ 8709] = 174;
assign img[ 8710] = 138;
assign img[ 8711] = 136;
assign img[ 8712] = 168;
assign img[ 8713] = 170;
assign img[ 8714] = 186;
assign img[ 8715] = 153;
assign img[ 8716] = 153;
assign img[ 8717] = 153;
assign img[ 8718] = 137;
assign img[ 8719] = 138;
assign img[ 8720] = 136;
assign img[ 8721] = 154;
assign img[ 8722] = 136;
assign img[ 8723] = 250;
assign img[ 8724] = 127;
assign img[ 8725] = 255;
assign img[ 8726] = 221;
assign img[ 8727] = 221;
assign img[ 8728] = 221;
assign img[ 8729] = 253;
assign img[ 8730] = 191;
assign img[ 8731] = 153;
assign img[ 8732] = 153;
assign img[ 8733] = 153;
assign img[ 8734] = 185;
assign img[ 8735] = 171;
assign img[ 8736] = 186;
assign img[ 8737] = 187;
assign img[ 8738] = 251;
assign img[ 8739] = 255;
assign img[ 8740] = 255;
assign img[ 8741] = 254;
assign img[ 8742] = 254;
assign img[ 8743] = 255;
assign img[ 8744] = 255;
assign img[ 8745] = 255;
assign img[ 8746] = 223;
assign img[ 8747] = 255;
assign img[ 8748] = 255;
assign img[ 8749] = 255;
assign img[ 8750] = 153;
assign img[ 8751] = 255;
assign img[ 8752] = 255;
assign img[ 8753] = 175;
assign img[ 8754] = 186;
assign img[ 8755] = 187;
assign img[ 8756] = 155;
assign img[ 8757] = 221;
assign img[ 8758] = 253;
assign img[ 8759] = 255;
assign img[ 8760] = 255;
assign img[ 8761] = 223;
assign img[ 8762] = 221;
assign img[ 8763] = 204;
assign img[ 8764] = 220;
assign img[ 8765] = 157;
assign img[ 8766] = 233;
assign img[ 8767] = 206;
assign img[ 8768] = 204;
assign img[ 8769] = 236;
assign img[ 8770] = 206;
assign img[ 8771] = 204;
assign img[ 8772] = 204;
assign img[ 8773] = 206;
assign img[ 8774] = 238;
assign img[ 8775] = 255;
assign img[ 8776] = 255;
assign img[ 8777] = 255;
assign img[ 8778] = 255;
assign img[ 8779] = 238;
assign img[ 8780] = 238;
assign img[ 8781] = 174;
assign img[ 8782] = 170;
assign img[ 8783] = 170;
assign img[ 8784] = 170;
assign img[ 8785] = 170;
assign img[ 8786] = 170;
assign img[ 8787] = 171;
assign img[ 8788] = 187;
assign img[ 8789] = 187;
assign img[ 8790] = 251;
assign img[ 8791] = 255;
assign img[ 8792] = 255;
assign img[ 8793] = 255;
assign img[ 8794] = 255;
assign img[ 8795] = 239;
assign img[ 8796] = 238;
assign img[ 8797] = 254;
assign img[ 8798] = 191;
assign img[ 8799] = 187;
assign img[ 8800] = 187;
assign img[ 8801] = 171;
assign img[ 8802] = 170;
assign img[ 8803] = 170;
assign img[ 8804] = 138;
assign img[ 8805] = 138;
assign img[ 8806] = 186;
assign img[ 8807] = 155;
assign img[ 8808] = 201;
assign img[ 8809] = 207;
assign img[ 8810] = 136;
assign img[ 8811] = 156;
assign img[ 8812] = 252;
assign img[ 8813] = 255;
assign img[ 8814] = 187;
assign img[ 8815] = 187;
assign img[ 8816] = 136;
assign img[ 8817] = 136;
assign img[ 8818] = 136;
assign img[ 8819] = 136;
assign img[ 8820] = 136;
assign img[ 8821] = 152;
assign img[ 8822] = 153;
assign img[ 8823] = 185;
assign img[ 8824] = 155;
assign img[ 8825] = 153;
assign img[ 8826] = 185;
assign img[ 8827] = 187;
assign img[ 8828] = 187;
assign img[ 8829] = 191;
assign img[ 8830] = 223;
assign img[ 8831] = 255;
assign img[ 8832] = 96;
assign img[ 8833] = 255;
assign img[ 8834] = 255;
assign img[ 8835] = 223;
assign img[ 8836] = 205;
assign img[ 8837] = 156;
assign img[ 8838] = 251;
assign img[ 8839] = 175;
assign img[ 8840] = 250;
assign img[ 8841] = 223;
assign img[ 8842] = 253;
assign img[ 8843] = 191;
assign img[ 8844] = 170;
assign img[ 8845] = 187;
assign img[ 8846] = 155;
assign img[ 8847] = 153;
assign img[ 8848] = 153;
assign img[ 8849] = 153;
assign img[ 8850] = 217;
assign img[ 8851] = 157;
assign img[ 8852] = 136;
assign img[ 8853] = 217;
assign img[ 8854] = 185;
assign img[ 8855] = 187;
assign img[ 8856] = 187;
assign img[ 8857] = 251;
assign img[ 8858] = 27;
assign img[ 8859] = 1;
assign img[ 8860] = 160;
assign img[ 8861] = 170;
assign img[ 8862] = 154;
assign img[ 8863] = 153;
assign img[ 8864] = 49;
assign img[ 8865] = 3;
assign img[ 8866] = 0;
assign img[ 8867] = 238;
assign img[ 8868] = 238;
assign img[ 8869] = 238;
assign img[ 8870] = 238;
assign img[ 8871] = 238;
assign img[ 8872] = 238;
assign img[ 8873] = 238;
assign img[ 8874] = 255;
assign img[ 8875] = 255;
assign img[ 8876] = 239;
assign img[ 8877] = 138;
assign img[ 8878] = 170;
assign img[ 8879] = 171;
assign img[ 8880] = 187;
assign img[ 8881] = 187;
assign img[ 8882] = 155;
assign img[ 8883] = 221;
assign img[ 8884] = 141;
assign img[ 8885] = 238;
assign img[ 8886] = 238;
assign img[ 8887] = 238;
assign img[ 8888] = 238;
assign img[ 8889] = 238;
assign img[ 8890] = 206;
assign img[ 8891] = 221;
assign img[ 8892] = 221;
assign img[ 8893] = 141;
assign img[ 8894] = 136;
assign img[ 8895] = 153;
assign img[ 8896] = 185;
assign img[ 8897] = 187;
assign img[ 8898] = 153;
assign img[ 8899] = 217;
assign img[ 8900] = 221;
assign img[ 8901] = 221;
assign img[ 8902] = 253;
assign img[ 8903] = 255;
assign img[ 8904] = 238;
assign img[ 8905] = 255;
assign img[ 8906] = 255;
assign img[ 8907] = 255;
assign img[ 8908] = 223;
assign img[ 8909] = 221;
assign img[ 8910] = 157;
assign img[ 8911] = 153;
assign img[ 8912] = 153;
assign img[ 8913] = 153;
assign img[ 8914] = 153;
assign img[ 8915] = 153;
assign img[ 8916] = 136;
assign img[ 8917] = 236;
assign img[ 8918] = 238;
assign img[ 8919] = 238;
assign img[ 8920] = 254;
assign img[ 8921] = 255;
assign img[ 8922] = 255;
assign img[ 8923] = 255;
assign img[ 8924] = 238;
assign img[ 8925] = 175;
assign img[ 8926] = 138;
assign img[ 8927] = 204;
assign img[ 8928] = 76;
assign img[ 8929] = 20;
assign img[ 8930] = 0;
assign img[ 8931] = 170;
assign img[ 8932] = 138;
assign img[ 8933] = 252;
assign img[ 8934] = 255;
assign img[ 8935] = 191;
assign img[ 8936] = 187;
assign img[ 8937] = 171;
assign img[ 8938] = 234;
assign img[ 8939] = 254;
assign img[ 8940] = 159;
assign img[ 8941] = 205;
assign img[ 8942] = 204;
assign img[ 8943] = 140;
assign img[ 8944] = 136;
assign img[ 8945] = 136;
assign img[ 8946] = 136;
assign img[ 8947] = 153;
assign img[ 8948] = 137;
assign img[ 8949] = 152;
assign img[ 8950] = 153;
assign img[ 8951] = 153;
assign img[ 8952] = 153;
assign img[ 8953] = 217;
assign img[ 8954] = 25;
assign img[ 8955] = 153;
assign img[ 8956] = 153;
assign img[ 8957] = 249;
assign img[ 8958] = 255;
assign img[ 8959] = 255;
assign img[ 8960] = 0;
assign img[ 8961] = 136;
assign img[ 8962] = 152;
assign img[ 8963] = 137;
assign img[ 8964] = 152;
assign img[ 8965] = 249;
assign img[ 8966] = 255;
assign img[ 8967] = 255;
assign img[ 8968] = 187;
assign img[ 8969] = 223;
assign img[ 8970] = 221;
assign img[ 8971] = 157;
assign img[ 8972] = 136;
assign img[ 8973] = 170;
assign img[ 8974] = 170;
assign img[ 8975] = 138;
assign img[ 8976] = 136;
assign img[ 8977] = 170;
assign img[ 8978] = 170;
assign img[ 8979] = 138;
assign img[ 8980] = 152;
assign img[ 8981] = 185;
assign img[ 8982] = 187;
assign img[ 8983] = 187;
assign img[ 8984] = 200;
assign img[ 8985] = 220;
assign img[ 8986] = 220;
assign img[ 8987] = 221;
assign img[ 8988] = 189;
assign img[ 8989] = 155;
assign img[ 8990] = 153;
assign img[ 8991] = 217;
assign img[ 8992] = 85;
assign img[ 8993] = 103;
assign img[ 8994] = 68;
assign img[ 8995] = 213;
assign img[ 8996] = 17;
assign img[ 8997] = 251;
assign img[ 8998] = 187;
assign img[ 8999] = 187;
assign img[ 9000] = 251;
assign img[ 9001] = 255;
assign img[ 9002] = 223;
assign img[ 9003] = 255;
assign img[ 9004] = 255;
assign img[ 9005] = 255;
assign img[ 9006] = 205;
assign img[ 9007] = 253;
assign img[ 9008] = 223;
assign img[ 9009] = 253;
assign img[ 9010] = 223;
assign img[ 9011] = 237;
assign img[ 9012] = 204;
assign img[ 9013] = 236;
assign img[ 9014] = 238;
assign img[ 9015] = 238;
assign img[ 9016] = 238;
assign img[ 9017] = 255;
assign img[ 9018] = 206;
assign img[ 9019] = 204;
assign img[ 9020] = 236;
assign img[ 9021] = 174;
assign img[ 9022] = 136;
assign img[ 9023] = 136;
assign img[ 9024] = 216;
assign img[ 9025] = 173;
assign img[ 9026] = 170;
assign img[ 9027] = 234;
assign img[ 9028] = 234;
assign img[ 9029] = 206;
assign img[ 9030] = 204;
assign img[ 9031] = 204;
assign img[ 9032] = 238;
assign img[ 9033] = 238;
assign img[ 9034] = 238;
assign img[ 9035] = 207;
assign img[ 9036] = 220;
assign img[ 9037] = 221;
assign img[ 9038] = 185;
assign img[ 9039] = 187;
assign img[ 9040] = 187;
assign img[ 9041] = 187;
assign img[ 9042] = 136;
assign img[ 9043] = 136;
assign img[ 9044] = 168;
assign img[ 9045] = 138;
assign img[ 9046] = 236;
assign img[ 9047] = 238;
assign img[ 9048] = 174;
assign img[ 9049] = 170;
assign img[ 9050] = 186;
assign img[ 9051] = 155;
assign img[ 9052] = 153;
assign img[ 9053] = 187;
assign img[ 9054] = 235;
assign img[ 9055] = 255;
assign img[ 9056] = 127;
assign img[ 9057] = 135;
assign img[ 9058] = 128;
assign img[ 9059] = 168;
assign img[ 9060] = 170;
assign img[ 9061] = 186;
assign img[ 9062] = 251;
assign img[ 9063] = 223;
assign img[ 9064] = 204;
assign img[ 9065] = 140;
assign img[ 9066] = 184;
assign img[ 9067] = 155;
assign img[ 9068] = 136;
assign img[ 9069] = 136;
assign img[ 9070] = 136;
assign img[ 9071] = 136;
assign img[ 9072] = 136;
assign img[ 9073] = 168;
assign img[ 9074] = 170;
assign img[ 9075] = 152;
assign img[ 9076] = 137;
assign img[ 9077] = 152;
assign img[ 9078] = 153;
assign img[ 9079] = 217;
assign img[ 9080] = 221;
assign img[ 9081] = 221;
assign img[ 9082] = 93;
assign img[ 9083] = 21;
assign img[ 9084] = 1;
assign img[ 9085] = 136;
assign img[ 9086] = 136;
assign img[ 9087] = 236;
assign img[ 9088] = 96;
assign img[ 9089] = 238;
assign img[ 9090] = 186;
assign img[ 9091] = 139;
assign img[ 9092] = 136;
assign img[ 9093] = 136;
assign img[ 9094] = 248;
assign img[ 9095] = 255;
assign img[ 9096] = 137;
assign img[ 9097] = 170;
assign img[ 9098] = 154;
assign img[ 9099] = 153;
assign img[ 9100] = 153;
assign img[ 9101] = 137;
assign img[ 9102] = 136;
assign img[ 9103] = 137;
assign img[ 9104] = 136;
assign img[ 9105] = 136;
assign img[ 9106] = 168;
assign img[ 9107] = 170;
assign img[ 9108] = 136;
assign img[ 9109] = 136;
assign img[ 9110] = 152;
assign img[ 9111] = 185;
assign img[ 9112] = 187;
assign img[ 9113] = 251;
assign img[ 9114] = 93;
assign img[ 9115] = 85;
assign img[ 9116] = 100;
assign img[ 9117] = 179;
assign img[ 9118] = 19;
assign img[ 9119] = 251;
assign img[ 9120] = 255;
assign img[ 9121] = 95;
assign img[ 9122] = 81;
assign img[ 9123] = 221;
assign img[ 9124] = 204;
assign img[ 9125] = 238;
assign img[ 9126] = 238;
assign img[ 9127] = 255;
assign img[ 9128] = 255;
assign img[ 9129] = 255;
assign img[ 9130] = 255;
assign img[ 9131] = 239;
assign img[ 9132] = 154;
assign img[ 9133] = 137;
assign img[ 9134] = 216;
assign img[ 9135] = 221;
assign img[ 9136] = 153;
assign img[ 9137] = 219;
assign img[ 9138] = 200;
assign img[ 9139] = 204;
assign img[ 9140] = 220;
assign img[ 9141] = 221;
assign img[ 9142] = 221;
assign img[ 9143] = 255;
assign img[ 9144] = 255;
assign img[ 9145] = 255;
assign img[ 9146] = 255;
assign img[ 9147] = 255;
assign img[ 9148] = 223;
assign img[ 9149] = 221;
assign img[ 9150] = 187;
assign img[ 9151] = 187;
assign img[ 9152] = 187;
assign img[ 9153] = 191;
assign img[ 9154] = 139;
assign img[ 9155] = 136;
assign img[ 9156] = 168;
assign img[ 9157] = 255;
assign img[ 9158] = 255;
assign img[ 9159] = 239;
assign img[ 9160] = 238;
assign img[ 9161] = 238;
assign img[ 9162] = 238;
assign img[ 9163] = 238;
assign img[ 9164] = 238;
assign img[ 9165] = 206;
assign img[ 9166] = 204;
assign img[ 9167] = 254;
assign img[ 9168] = 239;
assign img[ 9169] = 238;
assign img[ 9170] = 141;
assign img[ 9171] = 153;
assign img[ 9172] = 153;
assign img[ 9173] = 170;
assign img[ 9174] = 234;
assign img[ 9175] = 238;
assign img[ 9176] = 238;
assign img[ 9177] = 238;
assign img[ 9178] = 222;
assign img[ 9179] = 255;
assign img[ 9180] = 238;
assign img[ 9181] = 190;
assign img[ 9182] = 170;
assign img[ 9183] = 255;
assign img[ 9184] = 255;
assign img[ 9185] = 191;
assign img[ 9186] = 153;
assign img[ 9187] = 157;
assign img[ 9188] = 137;
assign img[ 9189] = 136;
assign img[ 9190] = 236;
assign img[ 9191] = 174;
assign img[ 9192] = 170;
assign img[ 9193] = 170;
assign img[ 9194] = 152;
assign img[ 9195] = 187;
assign img[ 9196] = 137;
assign img[ 9197] = 136;
assign img[ 9198] = 152;
assign img[ 9199] = 137;
assign img[ 9200] = 136;
assign img[ 9201] = 152;
assign img[ 9202] = 153;
assign img[ 9203] = 136;
assign img[ 9204] = 136;
assign img[ 9205] = 136;
assign img[ 9206] = 136;
assign img[ 9207] = 136;
assign img[ 9208] = 152;
assign img[ 9209] = 253;
assign img[ 9210] = 191;
assign img[ 9211] = 155;
assign img[ 9212] = 153;
assign img[ 9213] = 185;
assign img[ 9214] = 187;
assign img[ 9215] = 251;
assign img[ 9216] = 16;
assign img[ 9217] = 3;
assign img[ 9218] = 0;
assign img[ 9219] = 138;
assign img[ 9220] = 184;
assign img[ 9221] = 155;
assign img[ 9222] = 89;
assign img[ 9223] = 213;
assign img[ 9224] = 185;
assign img[ 9225] = 175;
assign img[ 9226] = 186;
assign img[ 9227] = 137;
assign img[ 9228] = 136;
assign img[ 9229] = 136;
assign img[ 9230] = 136;
assign img[ 9231] = 136;
assign img[ 9232] = 136;
assign img[ 9233] = 138;
assign img[ 9234] = 136;
assign img[ 9235] = 136;
assign img[ 9236] = 152;
assign img[ 9237] = 153;
assign img[ 9238] = 153;
assign img[ 9239] = 153;
assign img[ 9240] = 169;
assign img[ 9241] = 234;
assign img[ 9242] = 94;
assign img[ 9243] = 85;
assign img[ 9244] = 85;
assign img[ 9245] = 213;
assign img[ 9246] = 213;
assign img[ 9247] = 221;
assign img[ 9248] = 236;
assign img[ 9249] = 255;
assign img[ 9250] = 171;
assign img[ 9251] = 170;
assign img[ 9252] = 170;
assign img[ 9253] = 235;
assign img[ 9254] = 238;
assign img[ 9255] = 238;
assign img[ 9256] = 238;
assign img[ 9257] = 238;
assign img[ 9258] = 238;
assign img[ 9259] = 238;
assign img[ 9260] = 138;
assign img[ 9261] = 136;
assign img[ 9262] = 216;
assign img[ 9263] = 221;
assign img[ 9264] = 236;
assign img[ 9265] = 255;
assign img[ 9266] = 223;
assign img[ 9267] = 189;
assign img[ 9268] = 187;
assign img[ 9269] = 255;
assign img[ 9270] = 254;
assign img[ 9271] = 255;
assign img[ 9272] = 254;
assign img[ 9273] = 254;
assign img[ 9274] = 254;
assign img[ 9275] = 255;
assign img[ 9276] = 221;
assign img[ 9277] = 141;
assign img[ 9278] = 204;
assign img[ 9279] = 200;
assign img[ 9280] = 200;
assign img[ 9281] = 204;
assign img[ 9282] = 136;
assign img[ 9283] = 200;
assign img[ 9284] = 220;
assign img[ 9285] = 189;
assign img[ 9286] = 187;
assign img[ 9287] = 255;
assign img[ 9288] = 255;
assign img[ 9289] = 255;
assign img[ 9290] = 255;
assign img[ 9291] = 207;
assign img[ 9292] = 238;
assign img[ 9293] = 159;
assign img[ 9294] = 221;
assign img[ 9295] = 255;
assign img[ 9296] = 239;
assign img[ 9297] = 206;
assign img[ 9298] = 140;
assign img[ 9299] = 142;
assign img[ 9300] = 186;
assign img[ 9301] = 251;
assign img[ 9302] = 255;
assign img[ 9303] = 255;
assign img[ 9304] = 239;
assign img[ 9305] = 238;
assign img[ 9306] = 238;
assign img[ 9307] = 190;
assign img[ 9308] = 187;
assign img[ 9309] = 187;
assign img[ 9310] = 138;
assign img[ 9311] = 186;
assign img[ 9312] = 234;
assign img[ 9313] = 142;
assign img[ 9314] = 136;
assign img[ 9315] = 152;
assign img[ 9316] = 137;
assign img[ 9317] = 136;
assign img[ 9318] = 204;
assign img[ 9319] = 239;
assign img[ 9320] = 170;
assign img[ 9321] = 170;
assign img[ 9322] = 186;
assign img[ 9323] = 187;
assign img[ 9324] = 137;
assign img[ 9325] = 136;
assign img[ 9326] = 136;
assign img[ 9327] = 137;
assign img[ 9328] = 152;
assign img[ 9329] = 153;
assign img[ 9330] = 249;
assign img[ 9331] = 255;
assign img[ 9332] = 191;
assign img[ 9333] = 187;
assign img[ 9334] = 153;
assign img[ 9335] = 185;
assign img[ 9336] = 155;
assign img[ 9337] = 185;
assign img[ 9338] = 59;
assign img[ 9339] = 35;
assign img[ 9340] = 0;
assign img[ 9341] = 152;
assign img[ 9342] = 153;
assign img[ 9343] = 185;
assign img[ 9344] = 0;
assign img[ 9345] = 204;
assign img[ 9346] = 140;
assign img[ 9347] = 136;
assign img[ 9348] = 136;
assign img[ 9349] = 152;
assign img[ 9350] = 153;
assign img[ 9351] = 153;
assign img[ 9352] = 200;
assign img[ 9353] = 140;
assign img[ 9354] = 153;
assign img[ 9355] = 153;
assign img[ 9356] = 136;
assign img[ 9357] = 136;
assign img[ 9358] = 168;
assign img[ 9359] = 138;
assign img[ 9360] = 136;
assign img[ 9361] = 136;
assign img[ 9362] = 184;
assign img[ 9363] = 187;
assign img[ 9364] = 170;
assign img[ 9365] = 170;
assign img[ 9366] = 170;
assign img[ 9367] = 170;
assign img[ 9368] = 170;
assign img[ 9369] = 186;
assign img[ 9370] = 171;
assign img[ 9371] = 138;
assign img[ 9372] = 152;
assign img[ 9373] = 187;
assign img[ 9374] = 155;
assign img[ 9375] = 221;
assign img[ 9376] = 76;
assign img[ 9377] = 204;
assign img[ 9378] = 220;
assign img[ 9379] = 185;
assign img[ 9380] = 187;
assign img[ 9381] = 171;
assign img[ 9382] = 234;
assign img[ 9383] = 206;
assign img[ 9384] = 236;
assign img[ 9385] = 206;
assign img[ 9386] = 236;
assign img[ 9387] = 174;
assign img[ 9388] = 170;
assign img[ 9389] = 154;
assign img[ 9390] = 201;
assign img[ 9391] = 254;
assign img[ 9392] = 223;
assign img[ 9393] = 253;
assign img[ 9394] = 171;
assign img[ 9395] = 170;
assign img[ 9396] = 234;
assign img[ 9397] = 238;
assign img[ 9398] = 238;
assign img[ 9399] = 238;
assign img[ 9400] = 206;
assign img[ 9401] = 255;
assign img[ 9402] = 255;
assign img[ 9403] = 191;
assign img[ 9404] = 153;
assign img[ 9405] = 157;
assign img[ 9406] = 221;
assign img[ 9407] = 205;
assign img[ 9408] = 221;
assign img[ 9409] = 140;
assign img[ 9410] = 136;
assign img[ 9411] = 136;
assign img[ 9412] = 136;
assign img[ 9413] = 185;
assign img[ 9414] = 219;
assign img[ 9415] = 205;
assign img[ 9416] = 236;
assign img[ 9417] = 255;
assign img[ 9418] = 255;
assign img[ 9419] = 255;
assign img[ 9420] = 205;
assign img[ 9421] = 187;
assign img[ 9422] = 221;
assign img[ 9423] = 221;
assign img[ 9424] = 153;
assign img[ 9425] = 185;
assign img[ 9426] = 170;
assign img[ 9427] = 171;
assign img[ 9428] = 187;
assign img[ 9429] = 171;
assign img[ 9430] = 186;
assign img[ 9431] = 255;
assign img[ 9432] = 255;
assign img[ 9433] = 255;
assign img[ 9434] = 255;
assign img[ 9435] = 255;
assign img[ 9436] = 255;
assign img[ 9437] = 223;
assign img[ 9438] = 153;
assign img[ 9439] = 221;
assign img[ 9440] = 205;
assign img[ 9441] = 206;
assign img[ 9442] = 136;
assign img[ 9443] = 136;
assign img[ 9444] = 136;
assign img[ 9445] = 140;
assign img[ 9446] = 168;
assign img[ 9447] = 171;
assign img[ 9448] = 187;
assign img[ 9449] = 171;
assign img[ 9450] = 187;
assign img[ 9451] = 155;
assign img[ 9452] = 139;
assign img[ 9453] = 136;
assign img[ 9454] = 136;
assign img[ 9455] = 136;
assign img[ 9456] = 136;
assign img[ 9457] = 136;
assign img[ 9458] = 136;
assign img[ 9459] = 136;
assign img[ 9460] = 136;
assign img[ 9461] = 136;
assign img[ 9462] = 152;
assign img[ 9463] = 221;
assign img[ 9464] = 221;
assign img[ 9465] = 221;
assign img[ 9466] = 136;
assign img[ 9467] = 136;
assign img[ 9468] = 136;
assign img[ 9469] = 168;
assign img[ 9470] = 170;
assign img[ 9471] = 250;
assign img[ 9472] = 0;
assign img[ 9473] = 155;
assign img[ 9474] = 153;
assign img[ 9475] = 155;
assign img[ 9476] = 185;
assign img[ 9477] = 155;
assign img[ 9478] = 217;
assign img[ 9479] = 221;
assign img[ 9480] = 185;
assign img[ 9481] = 223;
assign img[ 9482] = 157;
assign img[ 9483] = 137;
assign img[ 9484] = 136;
assign img[ 9485] = 168;
assign img[ 9486] = 170;
assign img[ 9487] = 136;
assign img[ 9488] = 200;
assign img[ 9489] = 204;
assign img[ 9490] = 236;
assign img[ 9491] = 142;
assign img[ 9492] = 136;
assign img[ 9493] = 136;
assign img[ 9494] = 152;
assign img[ 9495] = 185;
assign img[ 9496] = 155;
assign img[ 9497] = 153;
assign img[ 9498] = 153;
assign img[ 9499] = 153;
assign img[ 9500] = 185;
assign img[ 9501] = 139;
assign img[ 9502] = 136;
assign img[ 9503] = 200;
assign img[ 9504] = 212;
assign img[ 9505] = 221;
assign img[ 9506] = 221;
assign img[ 9507] = 157;
assign img[ 9508] = 153;
assign img[ 9509] = 191;
assign img[ 9510] = 187;
assign img[ 9511] = 255;
assign img[ 9512] = 255;
assign img[ 9513] = 255;
assign img[ 9514] = 191;
assign img[ 9515] = 187;
assign img[ 9516] = 187;
assign img[ 9517] = 153;
assign img[ 9518] = 233;
assign img[ 9519] = 206;
assign img[ 9520] = 236;
assign img[ 9521] = 175;
assign img[ 9522] = 171;
assign img[ 9523] = 170;
assign img[ 9524] = 136;
assign img[ 9525] = 234;
assign img[ 9526] = 238;
assign img[ 9527] = 238;
assign img[ 9528] = 206;
assign img[ 9529] = 204;
assign img[ 9530] = 136;
assign img[ 9531] = 136;
assign img[ 9532] = 136;
assign img[ 9533] = 140;
assign img[ 9534] = 136;
assign img[ 9535] = 232;
assign img[ 9536] = 238;
assign img[ 9537] = 206;
assign img[ 9538] = 204;
assign img[ 9539] = 136;
assign img[ 9540] = 136;
assign img[ 9541] = 137;
assign img[ 9542] = 153;
assign img[ 9543] = 217;
assign img[ 9544] = 253;
assign img[ 9545] = 255;
assign img[ 9546] = 239;
assign img[ 9547] = 238;
assign img[ 9548] = 186;
assign img[ 9549] = 171;
assign img[ 9550] = 170;
assign img[ 9551] = 234;
assign img[ 9552] = 254;
assign img[ 9553] = 255;
assign img[ 9554] = 174;
assign img[ 9555] = 170;
assign img[ 9556] = 170;
assign img[ 9557] = 170;
assign img[ 9558] = 234;
assign img[ 9559] = 238;
assign img[ 9560] = 238;
assign img[ 9561] = 238;
assign img[ 9562] = 238;
assign img[ 9563] = 206;
assign img[ 9564] = 156;
assign img[ 9565] = 155;
assign img[ 9566] = 169;
assign img[ 9567] = 238;
assign img[ 9568] = 126;
assign img[ 9569] = 247;
assign img[ 9570] = 153;
assign img[ 9571] = 253;
assign img[ 9572] = 155;
assign img[ 9573] = 153;
assign img[ 9574] = 153;
assign img[ 9575] = 136;
assign img[ 9576] = 168;
assign img[ 9577] = 170;
assign img[ 9578] = 152;
assign img[ 9579] = 153;
assign img[ 9580] = 249;
assign img[ 9581] = 255;
assign img[ 9582] = 155;
assign img[ 9583] = 217;
assign img[ 9584] = 255;
assign img[ 9585] = 191;
assign img[ 9586] = 255;
assign img[ 9587] = 191;
assign img[ 9588] = 153;
assign img[ 9589] = 153;
assign img[ 9590] = 153;
assign img[ 9591] = 205;
assign img[ 9592] = 204;
assign img[ 9593] = 253;
assign img[ 9594] = 191;
assign img[ 9595] = 139;
assign img[ 9596] = 136;
assign img[ 9597] = 168;
assign img[ 9598] = 138;
assign img[ 9599] = 186;
assign img[ 9600] = 0;
assign img[ 9601] = 136;
assign img[ 9602] = 136;
assign img[ 9603] = 136;
assign img[ 9604] = 136;
assign img[ 9605] = 136;
assign img[ 9606] = 152;
assign img[ 9607] = 159;
assign img[ 9608] = 153;
assign img[ 9609] = 187;
assign img[ 9610] = 155;
assign img[ 9611] = 153;
assign img[ 9612] = 136;
assign img[ 9613] = 153;
assign img[ 9614] = 168;
assign img[ 9615] = 139;
assign img[ 9616] = 136;
assign img[ 9617] = 170;
assign img[ 9618] = 186;
assign img[ 9619] = 155;
assign img[ 9620] = 153;
assign img[ 9621] = 200;
assign img[ 9622] = 136;
assign img[ 9623] = 186;
assign img[ 9624] = 171;
assign img[ 9625] = 186;
assign img[ 9626] = 27;
assign img[ 9627] = 0;
assign img[ 9628] = 186;
assign img[ 9629] = 187;
assign img[ 9630] = 171;
assign img[ 9631] = 186;
assign img[ 9632] = 243;
assign img[ 9633] = 255;
assign img[ 9634] = 191;
assign img[ 9635] = 187;
assign img[ 9636] = 155;
assign img[ 9637] = 153;
assign img[ 9638] = 249;
assign img[ 9639] = 255;
assign img[ 9640] = 255;
assign img[ 9641] = 255;
assign img[ 9642] = 223;
assign img[ 9643] = 141;
assign img[ 9644] = 136;
assign img[ 9645] = 172;
assign img[ 9646] = 170;
assign img[ 9647] = 152;
assign img[ 9648] = 217;
assign img[ 9649] = 221;
assign img[ 9650] = 204;
assign img[ 9651] = 136;
assign img[ 9652] = 136;
assign img[ 9653] = 236;
assign img[ 9654] = 254;
assign img[ 9655] = 255;
assign img[ 9656] = 255;
assign img[ 9657] = 255;
assign img[ 9658] = 159;
assign img[ 9659] = 171;
assign img[ 9660] = 234;
assign img[ 9661] = 190;
assign img[ 9662] = 171;
assign img[ 9663] = 238;
assign img[ 9664] = 238;
assign img[ 9665] = 238;
assign img[ 9666] = 206;
assign img[ 9667] = 204;
assign img[ 9668] = 156;
assign img[ 9669] = 153;
assign img[ 9670] = 249;
assign img[ 9671] = 223;
assign img[ 9672] = 253;
assign img[ 9673] = 255;
assign img[ 9674] = 255;
assign img[ 9675] = 255;
assign img[ 9676] = 157;
assign img[ 9677] = 185;
assign img[ 9678] = 187;
assign img[ 9679] = 251;
assign img[ 9680] = 153;
assign img[ 9681] = 137;
assign img[ 9682] = 136;
assign img[ 9683] = 138;
assign img[ 9684] = 136;
assign img[ 9685] = 136;
assign img[ 9686] = 232;
assign img[ 9687] = 238;
assign img[ 9688] = 222;
assign img[ 9689] = 255;
assign img[ 9690] = 223;
assign img[ 9691] = 157;
assign img[ 9692] = 253;
assign img[ 9693] = 191;
assign img[ 9694] = 187;
assign img[ 9695] = 137;
assign img[ 9696] = 136;
assign img[ 9697] = 1;
assign img[ 9698] = 49;
assign img[ 9699] = 187;
assign img[ 9700] = 155;
assign img[ 9701] = 137;
assign img[ 9702] = 184;
assign img[ 9703] = 187;
assign img[ 9704] = 139;
assign img[ 9705] = 136;
assign img[ 9706] = 217;
assign img[ 9707] = 172;
assign img[ 9708] = 136;
assign img[ 9709] = 152;
assign img[ 9710] = 153;
assign img[ 9711] = 153;
assign img[ 9712] = 153;
assign img[ 9713] = 185;
assign img[ 9714] = 171;
assign img[ 9715] = 154;
assign img[ 9716] = 137;
assign img[ 9717] = 140;
assign img[ 9718] = 168;
assign img[ 9719] = 202;
assign img[ 9720] = 220;
assign img[ 9721] = 253;
assign img[ 9722] = 59;
assign img[ 9723] = 187;
assign img[ 9724] = 136;
assign img[ 9725] = 170;
assign img[ 9726] = 170;
assign img[ 9727] = 154;
assign img[ 9728] = 0;
assign img[ 9729] = 241;
assign img[ 9730] = 255;
assign img[ 9731] = 255;
assign img[ 9732] = 170;
assign img[ 9733] = 186;
assign img[ 9734] = 153;
assign img[ 9735] = 169;
assign img[ 9736] = 234;
assign img[ 9737] = 239;
assign img[ 9738] = 170;
assign img[ 9739] = 139;
assign img[ 9740] = 153;
assign img[ 9741] = 169;
assign img[ 9742] = 170;
assign img[ 9743] = 138;
assign img[ 9744] = 136;
assign img[ 9745] = 170;
assign img[ 9746] = 170;
assign img[ 9747] = 250;
assign img[ 9748] = 187;
assign img[ 9749] = 187;
assign img[ 9750] = 187;
assign img[ 9751] = 251;
assign img[ 9752] = 140;
assign img[ 9753] = 238;
assign img[ 9754] = 238;
assign img[ 9755] = 254;
assign img[ 9756] = 137;
assign img[ 9757] = 153;
assign img[ 9758] = 136;
assign img[ 9759] = 236;
assign img[ 9760] = 76;
assign img[ 9761] = 236;
assign img[ 9762] = 238;
assign img[ 9763] = 254;
assign img[ 9764] = 239;
assign img[ 9765] = 152;
assign img[ 9766] = 153;
assign img[ 9767] = 255;
assign img[ 9768] = 238;
assign img[ 9769] = 238;
assign img[ 9770] = 238;
assign img[ 9771] = 255;
assign img[ 9772] = 170;
assign img[ 9773] = 170;
assign img[ 9774] = 234;
assign img[ 9775] = 254;
assign img[ 9776] = 255;
assign img[ 9777] = 255;
assign img[ 9778] = 239;
assign img[ 9779] = 174;
assign img[ 9780] = 187;
assign img[ 9781] = 255;
assign img[ 9782] = 239;
assign img[ 9783] = 238;
assign img[ 9784] = 238;
assign img[ 9785] = 255;
assign img[ 9786] = 255;
assign img[ 9787] = 255;
assign img[ 9788] = 255;
assign img[ 9789] = 239;
assign img[ 9790] = 238;
assign img[ 9791] = 238;
assign img[ 9792] = 220;
assign img[ 9793] = 253;
assign img[ 9794] = 255;
assign img[ 9795] = 255;
assign img[ 9796] = 155;
assign img[ 9797] = 153;
assign img[ 9798] = 137;
assign img[ 9799] = 136;
assign img[ 9800] = 232;
assign img[ 9801] = 255;
assign img[ 9802] = 238;
assign img[ 9803] = 238;
assign img[ 9804] = 170;
assign img[ 9805] = 170;
assign img[ 9806] = 170;
assign img[ 9807] = 187;
assign img[ 9808] = 155;
assign img[ 9809] = 217;
assign img[ 9810] = 204;
assign img[ 9811] = 157;
assign img[ 9812] = 169;
assign img[ 9813] = 187;
assign img[ 9814] = 251;
assign img[ 9815] = 255;
assign img[ 9816] = 239;
assign img[ 9817] = 254;
assign img[ 9818] = 223;
assign img[ 9819] = 221;
assign img[ 9820] = 236;
assign img[ 9821] = 255;
assign img[ 9822] = 136;
assign img[ 9823] = 137;
assign img[ 9824] = 184;
assign img[ 9825] = 174;
assign img[ 9826] = 254;
assign img[ 9827] = 255;
assign img[ 9828] = 187;
assign img[ 9829] = 159;
assign img[ 9830] = 253;
assign img[ 9831] = 191;
assign img[ 9832] = 238;
assign img[ 9833] = 238;
assign img[ 9834] = 254;
assign img[ 9835] = 159;
assign img[ 9836] = 251;
assign img[ 9837] = 239;
assign img[ 9838] = 170;
assign img[ 9839] = 170;
assign img[ 9840] = 154;
assign img[ 9841] = 136;
assign img[ 9842] = 170;
assign img[ 9843] = 138;
assign img[ 9844] = 136;
assign img[ 9845] = 152;
assign img[ 9846] = 169;
assign img[ 9847] = 250;
assign img[ 9848] = 175;
assign img[ 9849] = 170;
assign img[ 9850] = 170;
assign img[ 9851] = 138;
assign img[ 9852] = 152;
assign img[ 9853] = 169;
assign img[ 9854] = 170;
assign img[ 9855] = 138;
assign img[ 9856] = 32;
assign img[ 9857] = 138;
assign img[ 9858] = 168;
assign img[ 9859] = 171;
assign img[ 9860] = 136;
assign img[ 9861] = 153;
assign img[ 9862] = 137;
assign img[ 9863] = 168;
assign img[ 9864] = 234;
assign img[ 9865] = 238;
assign img[ 9866] = 220;
assign img[ 9867] = 221;
assign img[ 9868] = 153;
assign img[ 9869] = 185;
assign img[ 9870] = 155;
assign img[ 9871] = 137;
assign img[ 9872] = 136;
assign img[ 9873] = 170;
assign img[ 9874] = 170;
assign img[ 9875] = 139;
assign img[ 9876] = 136;
assign img[ 9877] = 168;
assign img[ 9878] = 170;
assign img[ 9879] = 170;
assign img[ 9880] = 170;
assign img[ 9881] = 187;
assign img[ 9882] = 139;
assign img[ 9883] = 204;
assign img[ 9884] = 238;
assign img[ 9885] = 174;
assign img[ 9886] = 156;
assign img[ 9887] = 221;
assign img[ 9888] = 157;
assign img[ 9889] = 136;
assign img[ 9890] = 168;
assign img[ 9891] = 186;
assign img[ 9892] = 171;
assign img[ 9893] = 238;
assign img[ 9894] = 238;
assign img[ 9895] = 238;
assign img[ 9896] = 238;
assign img[ 9897] = 254;
assign img[ 9898] = 174;
assign img[ 9899] = 138;
assign img[ 9900] = 170;
assign img[ 9901] = 170;
assign img[ 9902] = 234;
assign img[ 9903] = 206;
assign img[ 9904] = 220;
assign img[ 9905] = 221;
assign img[ 9906] = 221;
assign img[ 9907] = 157;
assign img[ 9908] = 153;
assign img[ 9909] = 253;
assign img[ 9910] = 255;
assign img[ 9911] = 255;
assign img[ 9912] = 255;
assign img[ 9913] = 255;
assign img[ 9914] = 204;
assign img[ 9915] = 204;
assign img[ 9916] = 136;
assign img[ 9917] = 153;
assign img[ 9918] = 153;
assign img[ 9919] = 202;
assign img[ 9920] = 204;
assign img[ 9921] = 172;
assign img[ 9922] = 186;
assign img[ 9923] = 155;
assign img[ 9924] = 153;
assign img[ 9925] = 153;
assign img[ 9926] = 201;
assign img[ 9927] = 253;
assign img[ 9928] = 255;
assign img[ 9929] = 239;
assign img[ 9930] = 238;
assign img[ 9931] = 255;
assign img[ 9932] = 153;
assign img[ 9933] = 153;
assign img[ 9934] = 217;
assign img[ 9935] = 221;
assign img[ 9936] = 221;
assign img[ 9937] = 253;
assign img[ 9938] = 174;
assign img[ 9939] = 170;
assign img[ 9940] = 138;
assign img[ 9941] = 136;
assign img[ 9942] = 232;
assign img[ 9943] = 238;
assign img[ 9944] = 254;
assign img[ 9945] = 239;
assign img[ 9946] = 238;
assign img[ 9947] = 238;
assign img[ 9948] = 254;
assign img[ 9949] = 239;
assign img[ 9950] = 254;
assign img[ 9951] = 171;
assign img[ 9952] = 200;
assign img[ 9953] = 238;
assign img[ 9954] = 254;
assign img[ 9955] = 239;
assign img[ 9956] = 204;
assign img[ 9957] = 204;
assign img[ 9958] = 204;
assign img[ 9959] = 159;
assign img[ 9960] = 255;
assign img[ 9961] = 187;
assign img[ 9962] = 187;
assign img[ 9963] = 155;
assign img[ 9964] = 137;
assign img[ 9965] = 153;
assign img[ 9966] = 169;
assign img[ 9967] = 170;
assign img[ 9968] = 186;
assign img[ 9969] = 153;
assign img[ 9970] = 185;
assign img[ 9971] = 155;
assign img[ 9972] = 137;
assign img[ 9973] = 136;
assign img[ 9974] = 136;
assign img[ 9975] = 238;
assign img[ 9976] = 238;
assign img[ 9977] = 142;
assign img[ 9978] = 136;
assign img[ 9979] = 136;
assign img[ 9980] = 136;
assign img[ 9981] = 184;
assign img[ 9982] = 187;
assign img[ 9983] = 171;
assign img[ 9984] = 0;
assign img[ 9985] = 136;
assign img[ 9986] = 136;
assign img[ 9987] = 139;
assign img[ 9988] = 136;
assign img[ 9989] = 153;
assign img[ 9990] = 217;
assign img[ 9991] = 221;
assign img[ 9992] = 253;
assign img[ 9993] = 191;
assign img[ 9994] = 187;
assign img[ 9995] = 187;
assign img[ 9996] = 187;
assign img[ 9997] = 187;
assign img[ 9998] = 170;
assign img[ 9999] = 136;
assign img[10000] = 136;
assign img[10001] = 153;
assign img[10002] = 153;
assign img[10003] = 139;
assign img[10004] = 152;
assign img[10005] = 153;
assign img[10006] = 153;
assign img[10007] = 187;
assign img[10008] = 187;
assign img[10009] = 187;
assign img[10010] = 187;
assign img[10011] = 219;
assign img[10012] = 221;
assign img[10013] = 205;
assign img[10014] = 168;
assign img[10015] = 170;
assign img[10016] = 138;
assign img[10017] = 170;
assign img[10018] = 170;
assign img[10019] = 170;
assign img[10020] = 186;
assign img[10021] = 171;
assign img[10022] = 170;
assign img[10023] = 170;
assign img[10024] = 234;
assign img[10025] = 238;
assign img[10026] = 174;
assign img[10027] = 254;
assign img[10028] = 31;
assign img[10029] = 153;
assign img[10030] = 251;
assign img[10031] = 159;
assign img[10032] = 168;
assign img[10033] = 223;
assign img[10034] = 157;
assign img[10035] = 153;
assign img[10036] = 187;
assign img[10037] = 187;
assign img[10038] = 235;
assign img[10039] = 238;
assign img[10040] = 238;
assign img[10041] = 174;
assign img[10042] = 136;
assign img[10043] = 184;
assign img[10044] = 187;
assign img[10045] = 139;
assign img[10046] = 168;
assign img[10047] = 186;
assign img[10048] = 187;
assign img[10049] = 187;
assign img[10050] = 170;
assign img[10051] = 170;
assign img[10052] = 170;
assign img[10053] = 170;
assign img[10054] = 186;
assign img[10055] = 249;
assign img[10056] = 238;
assign img[10057] = 255;
assign img[10058] = 204;
assign img[10059] = 157;
assign img[10060] = 153;
assign img[10061] = 171;
assign img[10062] = 234;
assign img[10063] = 221;
assign img[10064] = 205;
assign img[10065] = 204;
assign img[10066] = 156;
assign img[10067] = 153;
assign img[10068] = 137;
assign img[10069] = 168;
assign img[10070] = 234;
assign img[10071] = 238;
assign img[10072] = 238;
assign img[10073] = 238;
assign img[10074] = 190;
assign img[10075] = 174;
assign img[10076] = 153;
assign img[10077] = 137;
assign img[10078] = 187;
assign img[10079] = 155;
assign img[10080] = 153;
assign img[10081] = 187;
assign img[10082] = 187;
assign img[10083] = 187;
assign img[10084] = 235;
assign img[10085] = 238;
assign img[10086] = 170;
assign img[10087] = 170;
assign img[10088] = 170;
assign img[10089] = 170;
assign img[10090] = 186;
assign img[10091] = 155;
assign img[10092] = 153;
assign img[10093] = 153;
assign img[10094] = 153;
assign img[10095] = 153;
assign img[10096] = 153;
assign img[10097] = 153;
assign img[10098] = 137;
assign img[10099] = 138;
assign img[10100] = 186;
assign img[10101] = 187;
assign img[10102] = 170;
assign img[10103] = 234;
assign img[10104] = 190;
assign img[10105] = 187;
assign img[10106] = 27;
assign img[10107] = 19;
assign img[10108] = 1;
assign img[10109] = 136;
assign img[10110] = 136;
assign img[10111] = 136;
assign img[10112] = 0;
assign img[10113] = 136;
assign img[10114] = 200;
assign img[10115] = 140;
assign img[10116] = 136;
assign img[10117] = 136;
assign img[10118] = 184;
assign img[10119] = 175;
assign img[10120] = 238;
assign img[10121] = 238;
assign img[10122] = 187;
assign img[10123] = 137;
assign img[10124] = 152;
assign img[10125] = 169;
assign img[10126] = 154;
assign img[10127] = 153;
assign img[10128] = 153;
assign img[10129] = 185;
assign img[10130] = 187;
assign img[10131] = 187;
assign img[10132] = 170;
assign img[10133] = 234;
assign img[10134] = 204;
assign img[10135] = 172;
assign img[10136] = 138;
assign img[10137] = 168;
assign img[10138] = 138;
assign img[10139] = 136;
assign img[10140] = 184;
assign img[10141] = 155;
assign img[10142] = 136;
assign img[10143] = 185;
assign img[10144] = 251;
assign img[10145] = 255;
assign img[10146] = 239;
assign img[10147] = 191;
assign img[10148] = 155;
assign img[10149] = 187;
assign img[10150] = 251;
assign img[10151] = 255;
assign img[10152] = 255;
assign img[10153] = 255;
assign img[10154] = 255;
assign img[10155] = 159;
assign img[10156] = 136;
assign img[10157] = 138;
assign img[10158] = 216;
assign img[10159] = 159;
assign img[10160] = 217;
assign img[10161] = 221;
assign img[10162] = 140;
assign img[10163] = 187;
assign img[10164] = 171;
assign img[10165] = 238;
assign img[10166] = 238;
assign img[10167] = 238;
assign img[10168] = 206;
assign img[10169] = 238;
assign img[10170] = 143;
assign img[10171] = 169;
assign img[10172] = 202;
assign img[10173] = 204;
assign img[10174] = 136;
assign img[10175] = 136;
assign img[10176] = 152;
assign img[10177] = 153;
assign img[10178] = 153;
assign img[10179] = 153;
assign img[10180] = 185;
assign img[10181] = 139;
assign img[10182] = 232;
assign img[10183] = 238;
assign img[10184] = 238;
assign img[10185] = 255;
assign img[10186] = 205;
assign img[10187] = 174;
assign img[10188] = 170;
assign img[10189] = 174;
assign img[10190] = 138;
assign img[10191] = 204;
assign img[10192] = 156;
assign img[10193] = 221;
assign img[10194] = 221;
assign img[10195] = 253;
assign img[10196] = 155;
assign img[10197] = 153;
assign img[10198] = 249;
assign img[10199] = 255;
assign img[10200] = 255;
assign img[10201] = 255;
assign img[10202] = 191;
assign img[10203] = 155;
assign img[10204] = 153;
assign img[10205] = 153;
assign img[10206] = 153;
assign img[10207] = 253;
assign img[10208] = 255;
assign img[10209] = 191;
assign img[10210] = 137;
assign img[10211] = 168;
assign img[10212] = 136;
assign img[10213] = 136;
assign img[10214] = 184;
assign img[10215] = 155;
assign img[10216] = 168;
assign img[10217] = 154;
assign img[10218] = 136;
assign img[10219] = 168;
assign img[10220] = 250;
assign img[10221] = 255;
assign img[10222] = 187;
assign img[10223] = 171;
assign img[10224] = 170;
assign img[10225] = 170;
assign img[10226] = 170;
assign img[10227] = 170;
assign img[10228] = 170;
assign img[10229] = 170;
assign img[10230] = 136;
assign img[10231] = 250;
assign img[10232] = 221;
assign img[10233] = 221;
assign img[10234] = 157;
assign img[10235] = 153;
assign img[10236] = 249;
assign img[10237] = 255;
assign img[10238] = 157;
assign img[10239] = 153;
assign img[10240] = 0;
assign img[10241] = 138;
assign img[10242] = 152;
assign img[10243] = 171;
assign img[10244] = 136;
assign img[10245] = 138;
assign img[10246] = 216;
assign img[10247] = 157;
assign img[10248] = 153;
assign img[10249] = 137;
assign img[10250] = 168;
assign img[10251] = 138;
assign img[10252] = 186;
assign img[10253] = 153;
assign img[10254] = 185;
assign img[10255] = 139;
assign img[10256] = 153;
assign img[10257] = 171;
assign img[10258] = 170;
assign img[10259] = 170;
assign img[10260] = 186;
assign img[10261] = 187;
assign img[10262] = 187;
assign img[10263] = 187;
assign img[10264] = 187;
assign img[10265] = 155;
assign img[10266] = 153;
assign img[10267] = 137;
assign img[10268] = 136;
assign img[10269] = 170;
assign img[10270] = 186;
assign img[10271] = 235;
assign img[10272] = 10;
assign img[10273] = 0;
assign img[10274] = 152;
assign img[10275] = 153;
assign img[10276] = 185;
assign img[10277] = 187;
assign img[10278] = 171;
assign img[10279] = 255;
assign img[10280] = 255;
assign img[10281] = 255;
assign img[10282] = 143;
assign img[10283] = 154;
assign img[10284] = 187;
assign img[10285] = 187;
assign img[10286] = 187;
assign img[10287] = 155;
assign img[10288] = 137;
assign img[10289] = 170;
assign img[10290] = 138;
assign img[10291] = 153;
assign img[10292] = 153;
assign img[10293] = 217;
assign img[10294] = 221;
assign img[10295] = 255;
assign img[10296] = 255;
assign img[10297] = 223;
assign img[10298] = 221;
assign img[10299] = 217;
assign img[10300] = 204;
assign img[10301] = 157;
assign img[10302] = 153;
assign img[10303] = 217;
assign img[10304] = 200;
assign img[10305] = 220;
assign img[10306] = 221;
assign img[10307] = 220;
assign img[10308] = 204;
assign img[10309] = 204;
assign img[10310] = 204;
assign img[10311] = 204;
assign img[10312] = 236;
assign img[10313] = 238;
assign img[10314] = 187;
assign img[10315] = 155;
assign img[10316] = 153;
assign img[10317] = 153;
assign img[10318] = 153;
assign img[10319] = 251;
assign img[10320] = 255;
assign img[10321] = 255;
assign img[10322] = 159;
assign img[10323] = 171;
assign img[10324] = 186;
assign img[10325] = 187;
assign img[10326] = 234;
assign img[10327] = 238;
assign img[10328] = 206;
assign img[10329] = 221;
assign img[10330] = 204;
assign img[10331] = 206;
assign img[10332] = 184;
assign img[10333] = 223;
assign img[10334] = 185;
assign img[10335] = 153;
assign img[10336] = 217;
assign img[10337] = 255;
assign img[10338] = 187;
assign img[10339] = 187;
assign img[10340] = 139;
assign img[10341] = 136;
assign img[10342] = 136;
assign img[10343] = 168;
assign img[10344] = 250;
assign img[10345] = 239;
assign img[10346] = 170;
assign img[10347] = 170;
assign img[10348] = 136;
assign img[10349] = 136;
assign img[10350] = 168;
assign img[10351] = 138;
assign img[10352] = 136;
assign img[10353] = 168;
assign img[10354] = 138;
assign img[10355] = 136;
assign img[10356] = 152;
assign img[10357] = 153;
assign img[10358] = 185;
assign img[10359] = 171;
assign img[10360] = 170;
assign img[10361] = 234;
assign img[10362] = 30;
assign img[10363] = 1;
assign img[10364] = 34;
assign img[10365] = 170;
assign img[10366] = 170;
assign img[10367] = 170;
assign img[10368] = 0;
assign img[10369] = 0;
assign img[10370] = 32;
assign img[10371] = 170;
assign img[10372] = 136;
assign img[10373] = 168;
assign img[10374] = 250;
assign img[10375] = 55;
assign img[10376] = 115;
assign img[10377] = 255;
assign img[10378] = 255;
assign img[10379] = 207;
assign img[10380] = 136;
assign img[10381] = 153;
assign img[10382] = 153;
assign img[10383] = 153;
assign img[10384] = 136;
assign img[10385] = 152;
assign img[10386] = 249;
assign img[10387] = 159;
assign img[10388] = 170;
assign img[10389] = 170;
assign img[10390] = 152;
assign img[10391] = 137;
assign img[10392] = 152;
assign img[10393] = 187;
assign img[10394] = 155;
assign img[10395] = 153;
assign img[10396] = 185;
assign img[10397] = 187;
assign img[10398] = 187;
assign img[10399] = 187;
assign img[10400] = 27;
assign img[10401] = 17;
assign img[10402] = 145;
assign img[10403] = 185;
assign img[10404] = 155;
assign img[10405] = 185;
assign img[10406] = 251;
assign img[10407] = 223;
assign img[10408] = 253;
assign img[10409] = 255;
assign img[10410] = 255;
assign img[10411] = 191;
assign img[10412] = 153;
assign img[10413] = 191;
assign img[10414] = 217;
assign img[10415] = 159;
assign img[10416] = 255;
assign img[10417] = 255;
assign img[10418] = 171;
assign img[10419] = 138;
assign img[10420] = 170;
assign img[10421] = 170;
assign img[10422] = 170;
assign img[10423] = 238;
assign img[10424] = 254;
assign img[10425] = 255;
assign img[10426] = 187;
assign img[10427] = 251;
assign img[10428] = 139;
assign img[10429] = 136;
assign img[10430] = 136;
assign img[10431] = 136;
assign img[10432] = 136;
assign img[10433] = 206;
assign img[10434] = 136;
assign img[10435] = 136;
assign img[10436] = 136;
assign img[10437] = 153;
assign img[10438] = 153;
assign img[10439] = 185;
assign img[10440] = 251;
assign img[10441] = 255;
assign img[10442] = 187;
assign img[10443] = 155;
assign img[10444] = 153;
assign img[10445] = 153;
assign img[10446] = 168;
assign img[10447] = 170;
assign img[10448] = 155;
assign img[10449] = 153;
assign img[10450] = 153;
assign img[10451] = 153;
assign img[10452] = 153;
assign img[10453] = 153;
assign img[10454] = 249;
assign img[10455] = 255;
assign img[10456] = 255;
assign img[10457] = 255;
assign img[10458] = 191;
assign img[10459] = 155;
assign img[10460] = 185;
assign img[10461] = 187;
assign img[10462] = 153;
assign img[10463] = 153;
assign img[10464] = 153;
assign img[10465] = 159;
assign img[10466] = 251;
assign img[10467] = 187;
assign img[10468] = 155;
assign img[10469] = 153;
assign img[10470] = 217;
assign img[10471] = 191;
assign img[10472] = 171;
assign img[10473] = 170;
assign img[10474] = 170;
assign img[10475] = 174;
assign img[10476] = 170;
assign img[10477] = 136;
assign img[10478] = 136;
assign img[10479] = 136;
assign img[10480] = 136;
assign img[10481] = 140;
assign img[10482] = 136;
assign img[10483] = 153;
assign img[10484] = 153;
assign img[10485] = 153;
assign img[10486] = 153;
assign img[10487] = 221;
assign img[10488] = 173;
assign img[10489] = 170;
assign img[10490] = 170;
assign img[10491] = 170;
assign img[10492] = 136;
assign img[10493] = 168;
assign img[10494] = 170;
assign img[10495] = 170;
assign img[10496] = 0;
assign img[10497] = 136;
assign img[10498] = 168;
assign img[10499] = 138;
assign img[10500] = 8;
assign img[10501] = 128;
assign img[10502] = 232;
assign img[10503] = 223;
assign img[10504] = 153;
assign img[10505] = 221;
assign img[10506] = 157;
assign img[10507] = 153;
assign img[10508] = 153;
assign img[10509] = 153;
assign img[10510] = 153;
assign img[10511] = 137;
assign img[10512] = 136;
assign img[10513] = 136;
assign img[10514] = 136;
assign img[10515] = 140;
assign img[10516] = 184;
assign img[10517] = 153;
assign img[10518] = 153;
assign img[10519] = 153;
assign img[10520] = 169;
assign img[10521] = 170;
assign img[10522] = 152;
assign img[10523] = 249;
assign img[10524] = 238;
assign img[10525] = 254;
assign img[10526] = 157;
assign img[10527] = 221;
assign img[10528] = 249;
assign img[10529] = 207;
assign img[10530] = 204;
assign img[10531] = 236;
assign img[10532] = 142;
assign img[10533] = 136;
assign img[10534] = 152;
assign img[10535] = 201;
assign img[10536] = 236;
assign img[10537] = 238;
assign img[10538] = 174;
assign img[10539] = 138;
assign img[10540] = 168;
assign img[10541] = 170;
assign img[10542] = 152;
assign img[10543] = 157;
assign img[10544] = 205;
assign img[10545] = 220;
assign img[10546] = 253;
assign img[10547] = 239;
assign img[10548] = 238;
assign img[10549] = 174;
assign img[10550] = 138;
assign img[10551] = 238;
assign img[10552] = 238;
assign img[10553] = 223;
assign img[10554] = 255;
assign img[10555] = 223;
assign img[10556] = 255;
assign img[10557] = 221;
assign img[10558] = 153;
assign img[10559] = 221;
assign img[10560] = 221;
assign img[10561] = 221;
assign img[10562] = 221;
assign img[10563] = 205;
assign img[10564] = 204;
assign img[10565] = 204;
assign img[10566] = 204;
assign img[10567] = 185;
assign img[10568] = 251;
assign img[10569] = 255;
assign img[10570] = 221;
assign img[10571] = 159;
assign img[10572] = 153;
assign img[10573] = 175;
assign img[10574] = 206;
assign img[10575] = 204;
assign img[10576] = 157;
assign img[10577] = 153;
assign img[10578] = 153;
assign img[10579] = 153;
assign img[10580] = 187;
assign img[10581] = 187;
assign img[10582] = 234;
assign img[10583] = 255;
assign img[10584] = 255;
assign img[10585] = 187;
assign img[10586] = 153;
assign img[10587] = 153;
assign img[10588] = 185;
assign img[10589] = 187;
assign img[10590] = 217;
assign img[10591] = 253;
assign img[10592] = 221;
assign img[10593] = 255;
assign img[10594] = 255;
assign img[10595] = 223;
assign img[10596] = 236;
assign img[10597] = 206;
assign img[10598] = 136;
assign img[10599] = 136;
assign img[10600] = 136;
assign img[10601] = 187;
assign img[10602] = 153;
assign img[10603] = 155;
assign img[10604] = 153;
assign img[10605] = 153;
assign img[10606] = 153;
assign img[10607] = 153;
assign img[10608] = 153;
assign img[10609] = 153;
assign img[10610] = 185;
assign img[10611] = 187;
assign img[10612] = 187;
assign img[10613] = 153;
assign img[10614] = 137;
assign img[10615] = 136;
assign img[10616] = 136;
assign img[10617] = 253;
assign img[10618] = 63;
assign img[10619] = 19;
assign img[10620] = 17;
assign img[10621] = 129;
assign img[10622] = 136;
assign img[10623] = 136;
assign img[10624] = 0;
assign img[10625] = 128;
assign img[10626] = 248;
assign img[10627] = 191;
assign img[10628] = 187;
assign img[10629] = 187;
assign img[10630] = 251;
assign img[10631] = 175;
assign img[10632] = 170;
assign img[10633] = 170;
assign img[10634] = 136;
assign img[10635] = 170;
assign img[10636] = 136;
assign img[10637] = 169;
assign img[10638] = 187;
assign img[10639] = 187;
assign img[10640] = 187;
assign img[10641] = 187;
assign img[10642] = 234;
assign img[10643] = 191;
assign img[10644] = 187;
assign img[10645] = 187;
assign img[10646] = 153;
assign img[10647] = 153;
assign img[10648] = 137;
assign img[10649] = 238;
assign img[10650] = 46;
assign img[10651] = 50;
assign img[10652] = 179;
assign img[10653] = 187;
assign img[10654] = 138;
assign img[10655] = 217;
assign img[10656] = 9;
assign img[10657] = 64;
assign img[10658] = 36;
assign img[10659] = 2;
assign img[10660] = 128;
assign img[10661] = 169;
assign img[10662] = 235;
assign img[10663] = 204;
assign img[10664] = 236;
assign img[10665] = 254;
assign img[10666] = 206;
assign img[10667] = 204;
assign img[10668] = 204;
assign img[10669] = 221;
assign img[10670] = 253;
assign img[10671] = 255;
assign img[10672] = 187;
assign img[10673] = 255;
assign img[10674] = 171;
assign img[10675] = 170;
assign img[10676] = 170;
assign img[10677] = 234;
assign img[10678] = 238;
assign img[10679] = 238;
assign img[10680] = 190;
assign img[10681] = 155;
assign img[10682] = 153;
assign img[10683] = 185;
assign img[10684] = 234;
assign img[10685] = 174;
assign img[10686] = 186;
assign img[10687] = 187;
assign img[10688] = 187;
assign img[10689] = 187;
assign img[10690] = 187;
assign img[10691] = 187;
assign img[10692] = 170;
assign img[10693] = 138;
assign img[10694] = 136;
assign img[10695] = 136;
assign img[10696] = 232;
assign img[10697] = 255;
assign img[10698] = 255;
assign img[10699] = 255;
assign img[10700] = 187;
assign img[10701] = 187;
assign img[10702] = 168;
assign img[10703] = 170;
assign img[10704] = 152;
assign img[10705] = 253;
assign img[10706] = 255;
assign img[10707] = 206;
assign img[10708] = 204;
assign img[10709] = 204;
assign img[10710] = 236;
assign img[10711] = 238;
assign img[10712] = 238;
assign img[10713] = 206;
assign img[10714] = 236;
assign img[10715] = 254;
assign img[10716] = 171;
assign img[10717] = 170;
assign img[10718] = 202;
assign img[10719] = 140;
assign img[10720] = 200;
assign img[10721] = 157;
assign img[10722] = 185;
assign img[10723] = 187;
assign img[10724] = 187;
assign img[10725] = 239;
assign img[10726] = 220;
assign img[10727] = 253;
assign img[10728] = 187;
assign img[10729] = 187;
assign img[10730] = 187;
assign img[10731] = 191;
assign img[10732] = 187;
assign img[10733] = 251;
assign img[10734] = 137;
assign img[10735] = 136;
assign img[10736] = 136;
assign img[10737] = 170;
assign img[10738] = 170;
assign img[10739] = 186;
assign img[10740] = 171;
assign img[10741] = 170;
assign img[10742] = 154;
assign img[10743] = 187;
assign img[10744] = 170;
assign img[10745] = 250;
assign img[10746] = 138;
assign img[10747] = 136;
assign img[10748] = 136;
assign img[10749] = 136;
assign img[10750] = 136;
assign img[10751] = 153;
assign img[10752] = 16;
assign img[10753] = 155;
assign img[10754] = 136;
assign img[10755] = 138;
assign img[10756] = 136;
assign img[10757] = 152;
assign img[10758] = 153;
assign img[10759] = 153;
assign img[10760] = 153;
assign img[10761] = 141;
assign img[10762] = 136;
assign img[10763] = 170;
assign img[10764] = 186;
assign img[10765] = 153;
assign img[10766] = 136;
assign img[10767] = 137;
assign img[10768] = 152;
assign img[10769] = 153;
assign img[10770] = 137;
assign img[10771] = 137;
assign img[10772] = 136;
assign img[10773] = 136;
assign img[10774] = 152;
assign img[10775] = 137;
assign img[10776] = 200;
assign img[10777] = 140;
assign img[10778] = 168;
assign img[10779] = 206;
assign img[10780] = 252;
assign img[10781] = 175;
assign img[10782] = 170;
assign img[10783] = 170;
assign img[10784] = 186;
assign img[10785] = 187;
assign img[10786] = 155;
assign img[10787] = 187;
assign img[10788] = 187;
assign img[10789] = 155;
assign img[10790] = 249;
assign img[10791] = 255;
assign img[10792] = 255;
assign img[10793] = 223;
assign img[10794] = 221;
assign img[10795] = 223;
assign img[10796] = 239;
assign img[10797] = 238;
assign img[10798] = 238;
assign img[10799] = 174;
assign img[10800] = 138;
assign img[10801] = 136;
assign img[10802] = 136;
assign img[10803] = 186;
assign img[10804] = 187;
assign img[10805] = 187;
assign img[10806] = 187;
assign img[10807] = 155;
assign img[10808] = 185;
assign img[10809] = 187;
assign img[10810] = 170;
assign img[10811] = 152;
assign img[10812] = 153;
assign img[10813] = 155;
assign img[10814] = 185;
assign img[10815] = 171;
assign img[10816] = 170;
assign img[10817] = 187;
assign img[10818] = 187;
assign img[10819] = 187;
assign img[10820] = 155;
assign img[10821] = 153;
assign img[10822] = 168;
assign img[10823] = 186;
assign img[10824] = 155;
assign img[10825] = 221;
assign img[10826] = 189;
assign img[10827] = 187;
assign img[10828] = 187;
assign img[10829] = 171;
assign img[10830] = 250;
assign img[10831] = 223;
assign img[10832] = 153;
assign img[10833] = 235;
assign img[10834] = 254;
assign img[10835] = 239;
assign img[10836] = 238;
assign img[10837] = 255;
assign img[10838] = 255;
assign img[10839] = 255;
assign img[10840] = 255;
assign img[10841] = 239;
assign img[10842] = 190;
assign img[10843] = 155;
assign img[10844] = 185;
assign img[10845] = 187;
assign img[10846] = 153;
assign img[10847] = 221;
assign img[10848] = 237;
assign img[10849] = 255;
assign img[10850] = 187;
assign img[10851] = 187;
assign img[10852] = 187;
assign img[10853] = 175;
assign img[10854] = 254;
assign img[10855] = 239;
assign img[10856] = 204;
assign img[10857] = 204;
assign img[10858] = 153;
assign img[10859] = 153;
assign img[10860] = 249;
assign img[10861] = 223;
assign img[10862] = 221;
assign img[10863] = 221;
assign img[10864] = 253;
assign img[10865] = 223;
assign img[10866] = 169;
assign img[10867] = 170;
assign img[10868] = 170;
assign img[10869] = 170;
assign img[10870] = 170;
assign img[10871] = 186;
assign img[10872] = 153;
assign img[10873] = 153;
assign img[10874] = 249;
assign img[10875] = 143;
assign img[10876] = 136;
assign img[10877] = 136;
assign img[10878] = 136;
assign img[10879] = 168;
assign img[10880] = 0;
assign img[10881] = 2;
assign img[10882] = 0;
assign img[10883] = 136;
assign img[10884] = 136;
assign img[10885] = 153;
assign img[10886] = 217;
assign img[10887] = 255;
assign img[10888] = 169;
assign img[10889] = 170;
assign img[10890] = 170;
assign img[10891] = 171;
assign img[10892] = 251;
assign img[10893] = 239;
assign img[10894] = 138;
assign img[10895] = 136;
assign img[10896] = 136;
assign img[10897] = 136;
assign img[10898] = 136;
assign img[10899] = 136;
assign img[10900] = 168;
assign img[10901] = 170;
assign img[10902] = 136;
assign img[10903] = 136;
assign img[10904] = 168;
assign img[10905] = 187;
assign img[10906] = 187;
assign img[10907] = 153;
assign img[10908] = 201;
assign img[10909] = 221;
assign img[10910] = 157;
assign img[10911] = 153;
assign img[10912] = 249;
assign img[10913] = 255;
assign img[10914] = 255;
assign img[10915] = 255;
assign img[10916] = 157;
assign img[10917] = 185;
assign img[10918] = 187;
assign img[10919] = 187;
assign img[10920] = 234;
assign img[10921] = 238;
assign img[10922] = 238;
assign img[10923] = 255;
assign img[10924] = 170;
assign img[10925] = 170;
assign img[10926] = 170;
assign img[10927] = 174;
assign img[10928] = 254;
assign img[10929] = 191;
assign img[10930] = 187;
assign img[10931] = 251;
assign img[10932] = 255;
assign img[10933] = 239;
assign img[10934] = 206;
assign img[10935] = 236;
assign img[10936] = 238;
assign img[10937] = 206;
assign img[10938] = 221;
assign img[10939] = 239;
assign img[10940] = 238;
assign img[10941] = 191;
assign img[10942] = 187;
assign img[10943] = 187;
assign img[10944] = 251;
assign img[10945] = 191;
assign img[10946] = 155;
assign img[10947] = 221;
assign img[10948] = 157;
assign img[10949] = 137;
assign img[10950] = 152;
assign img[10951] = 137;
assign img[10952] = 236;
assign img[10953] = 223;
assign img[10954] = 253;
assign img[10955] = 255;
assign img[10956] = 239;
assign img[10957] = 174;
assign img[10958] = 170;
assign img[10959] = 251;
assign img[10960] = 255;
assign img[10961] = 255;
assign img[10962] = 191;
assign img[10963] = 155;
assign img[10964] = 153;
assign img[10965] = 153;
assign img[10966] = 153;
assign img[10967] = 253;
assign img[10968] = 239;
assign img[10969] = 238;
assign img[10970] = 238;
assign img[10971] = 174;
assign img[10972] = 200;
assign img[10973] = 236;
assign img[10974] = 238;
assign img[10975] = 140;
assign img[10976] = 136;
assign img[10977] = 140;
assign img[10978] = 152;
assign img[10979] = 221;
assign img[10980] = 221;
assign img[10981] = 140;
assign img[10982] = 136;
assign img[10983] = 185;
assign img[10984] = 139;
assign img[10985] = 136;
assign img[10986] = 204;
assign img[10987] = 204;
assign img[10988] = 204;
assign img[10989] = 220;
assign img[10990] = 221;
assign img[10991] = 221;
assign img[10992] = 221;
assign img[10993] = 153;
assign img[10994] = 185;
assign img[10995] = 187;
assign img[10996] = 170;
assign img[10997] = 136;
assign img[10998] = 152;
assign img[10999] = 185;
assign img[11000] = 170;
assign img[11001] = 251;
assign img[11002] = 223;
assign img[11003] = 221;
assign img[11004] = 221;
assign img[11005] = 185;
assign img[11006] = 155;
assign img[11007] = 168;
assign img[11008] = 0;
assign img[11009] = 136;
assign img[11010] = 136;
assign img[11011] = 152;
assign img[11012] = 153;
assign img[11013] = 153;
assign img[11014] = 217;
assign img[11015] = 221;
assign img[11016] = 153;
assign img[11017] = 157;
assign img[11018] = 185;
assign img[11019] = 155;
assign img[11020] = 168;
assign img[11021] = 186;
assign img[11022] = 170;
assign img[11023] = 170;
assign img[11024] = 170;
assign img[11025] = 186;
assign img[11026] = 137;
assign img[11027] = 170;
assign img[11028] = 170;
assign img[11029] = 170;
assign img[11030] = 154;
assign img[11031] = 187;
assign img[11032] = 187;
assign img[11033] = 171;
assign img[11034] = 170;
assign img[11035] = 206;
assign img[11036] = 204;
assign img[11037] = 236;
assign img[11038] = 138;
assign img[11039] = 234;
assign img[11040] = 34;
assign img[11041] = 226;
assign img[11042] = 238;
assign img[11043] = 238;
assign img[11044] = 170;
assign img[11045] = 170;
assign img[11046] = 186;
assign img[11047] = 171;
assign img[11048] = 234;
assign img[11049] = 255;
assign img[11050] = 187;
assign img[11051] = 171;
assign img[11052] = 186;
assign img[11053] = 187;
assign img[11054] = 234;
assign img[11055] = 223;
assign img[11056] = 205;
assign img[11057] = 221;
assign img[11058] = 221;
assign img[11059] = 157;
assign img[11060] = 136;
assign img[11061] = 152;
assign img[11062] = 153;
assign img[11063] = 221;
assign img[11064] = 185;
assign img[11065] = 155;
assign img[11066] = 153;
assign img[11067] = 157;
assign img[11068] = 221;
assign img[11069] = 204;
assign img[11070] = 236;
assign img[11071] = 222;
assign img[11072] = 221;
assign img[11073] = 253;
assign img[11074] = 255;
assign img[11075] = 255;
assign img[11076] = 238;
assign img[11077] = 206;
assign img[11078] = 184;
assign img[11079] = 171;
assign img[11080] = 202;
assign img[11081] = 221;
assign img[11082] = 221;
assign img[11083] = 153;
assign img[11084] = 136;
assign img[11085] = 152;
assign img[11086] = 153;
assign img[11087] = 153;
assign img[11088] = 153;
assign img[11089] = 253;
assign img[11090] = 175;
assign img[11091] = 170;
assign img[11092] = 138;
assign img[11093] = 152;
assign img[11094] = 185;
assign img[11095] = 255;
assign img[11096] = 255;
assign img[11097] = 191;
assign img[11098] = 187;
assign img[11099] = 187;
assign img[11100] = 187;
assign img[11101] = 155;
assign img[11102] = 217;
assign img[11103] = 205;
assign img[11104] = 253;
assign img[11105] = 55;
assign img[11106] = 81;
assign img[11107] = 221;
assign img[11108] = 221;
assign img[11109] = 221;
assign img[11110] = 221;
assign img[11111] = 191;
assign img[11112] = 187;
assign img[11113] = 187;
assign img[11114] = 153;
assign img[11115] = 187;
assign img[11116] = 187;
assign img[11117] = 171;
assign img[11118] = 170;
assign img[11119] = 170;
assign img[11120] = 234;
assign img[11121] = 170;
assign img[11122] = 186;
assign img[11123] = 155;
assign img[11124] = 153;
assign img[11125] = 153;
assign img[11126] = 137;
assign img[11127] = 153;
assign img[11128] = 153;
assign img[11129] = 255;
assign img[11130] = 191;
assign img[11131] = 171;
assign img[11132] = 170;
assign img[11133] = 170;
assign img[11134] = 138;
assign img[11135] = 139;
assign img[11136] = 16;
assign img[11137] = 155;
assign img[11138] = 170;
assign img[11139] = 187;
assign img[11140] = 153;
assign img[11141] = 136;
assign img[11142] = 200;
assign img[11143] = 68;
assign img[11144] = 0;
assign img[11145] = 136;
assign img[11146] = 136;
assign img[11147] = 138;
assign img[11148] = 136;
assign img[11149] = 249;
assign img[11150] = 255;
assign img[11151] = 191;
assign img[11152] = 187;
assign img[11153] = 171;
assign img[11154] = 204;
assign img[11155] = 204;
assign img[11156] = 236;
assign img[11157] = 170;
assign img[11158] = 186;
assign img[11159] = 171;
assign img[11160] = 170;
assign img[11161] = 255;
assign img[11162] = 175;
assign img[11163] = 200;
assign img[11164] = 236;
assign img[11165] = 239;
assign img[11166] = 238;
assign img[11167] = 136;
assign img[11168] = 136;
assign img[11169] = 136;
assign img[11170] = 152;
assign img[11171] = 205;
assign img[11172] = 156;
assign img[11173] = 153;
assign img[11174] = 153;
assign img[11175] = 205;
assign img[11176] = 236;
assign img[11177] = 223;
assign img[11178] = 221;
assign img[11179] = 221;
assign img[11180] = 221;
assign img[11181] = 221;
assign img[11182] = 253;
assign img[11183] = 223;
assign img[11184] = 253;
assign img[11185] = 255;
assign img[11186] = 255;
assign img[11187] = 255;
assign img[11188] = 137;
assign img[11189] = 217;
assign img[11190] = 217;
assign img[11191] = 253;
assign img[11192] = 239;
assign img[11193] = 238;
assign img[11194] = 238;
assign img[11195] = 170;
assign img[11196] = 234;
assign img[11197] = 238;
assign img[11198] = 170;
assign img[11199] = 206;
assign img[11200] = 204;
assign img[11201] = 220;
assign img[11202] = 253;
assign img[11203] = 255;
assign img[11204] = 239;
assign img[11205] = 174;
assign img[11206] = 186;
assign img[11207] = 191;
assign img[11208] = 238;
assign img[11209] = 206;
assign img[11210] = 204;
assign img[11211] = 205;
assign img[11212] = 204;
assign img[11213] = 204;
assign img[11214] = 236;
assign img[11215] = 255;
assign img[11216] = 223;
assign img[11217] = 221;
assign img[11218] = 204;
assign img[11219] = 204;
assign img[11220] = 152;
assign img[11221] = 153;
assign img[11222] = 217;
assign img[11223] = 253;
assign img[11224] = 223;
assign img[11225] = 205;
assign img[11226] = 220;
assign img[11227] = 153;
assign img[11228] = 249;
assign img[11229] = 221;
assign img[11230] = 205;
assign img[11231] = 140;
assign img[11232] = 136;
assign img[11233] = 152;
assign img[11234] = 137;
assign img[11235] = 152;
assign img[11236] = 153;
assign img[11237] = 153;
assign img[11238] = 232;
assign img[11239] = 255;
assign img[11240] = 239;
assign img[11241] = 238;
assign img[11242] = 186;
assign img[11243] = 187;
assign img[11244] = 155;
assign img[11245] = 200;
assign img[11246] = 204;
assign img[11247] = 222;
assign img[11248] = 205;
assign img[11249] = 253;
assign img[11250] = 254;
assign img[11251] = 255;
assign img[11252] = 153;
assign img[11253] = 185;
assign img[11254] = 187;
assign img[11255] = 187;
assign img[11256] = 187;
assign img[11257] = 255;
assign img[11258] = 255;
assign img[11259] = 207;
assign img[11260] = 204;
assign img[11261] = 185;
assign img[11262] = 171;
assign img[11263] = 170;
assign img[11264] = 48;
assign img[11265] = 139;
assign img[11266] = 136;
assign img[11267] = 8;
assign img[11268] = 136;
assign img[11269] = 136;
assign img[11270] = 136;
assign img[11271] = 168;
assign img[11272] = 254;
assign img[11273] = 255;
assign img[11274] = 221;
assign img[11275] = 204;
assign img[11276] = 236;
assign img[11277] = 238;
assign img[11278] = 170;
assign img[11279] = 187;
assign img[11280] = 137;
assign img[11281] = 136;
assign img[11282] = 168;
assign img[11283] = 138;
assign img[11284] = 168;
assign img[11285] = 186;
assign img[11286] = 187;
assign img[11287] = 234;
assign img[11288] = 204;
assign img[11289] = 140;
assign img[11290] = 136;
assign img[11291] = 234;
assign img[11292] = 206;
assign img[11293] = 204;
assign img[11294] = 152;
assign img[11295] = 153;
assign img[11296] = 25;
assign img[11297] = 221;
assign img[11298] = 204;
assign img[11299] = 190;
assign img[11300] = 155;
assign img[11301] = 137;
assign img[11302] = 152;
assign img[11303] = 155;
assign img[11304] = 251;
assign img[11305] = 255;
assign img[11306] = 255;
assign img[11307] = 187;
assign img[11308] = 187;
assign img[11309] = 171;
assign img[11310] = 170;
assign img[11311] = 170;
assign img[11312] = 234;
assign img[11313] = 191;
assign img[11314] = 171;
assign img[11315] = 170;
assign img[11316] = 138;
assign img[11317] = 206;
assign img[11318] = 236;
assign img[11319] = 206;
assign img[11320] = 204;
assign img[11321] = 236;
assign img[11322] = 238;
assign img[11323] = 238;
assign img[11324] = 206;
assign img[11325] = 204;
assign img[11326] = 204;
assign img[11327] = 204;
assign img[11328] = 204;
assign img[11329] = 204;
assign img[11330] = 204;
assign img[11331] = 204;
assign img[11332] = 140;
assign img[11333] = 138;
assign img[11334] = 136;
assign img[11335] = 234;
assign img[11336] = 254;
assign img[11337] = 221;
assign img[11338] = 221;
assign img[11339] = 221;
assign img[11340] = 205;
assign img[11341] = 141;
assign img[11342] = 168;
assign img[11343] = 202;
assign img[11344] = 136;
assign img[11345] = 234;
assign img[11346] = 170;
assign img[11347] = 170;
assign img[11348] = 187;
assign img[11349] = 187;
assign img[11350] = 137;
assign img[11351] = 238;
assign img[11352] = 238;
assign img[11353] = 174;
assign img[11354] = 170;
assign img[11355] = 138;
assign img[11356] = 185;
assign img[11357] = 187;
assign img[11358] = 251;
assign img[11359] = 255;
assign img[11360] = 255;
assign img[11361] = 23;
assign img[11362] = 51;
assign img[11363] = 187;
assign img[11364] = 235;
assign img[11365] = 174;
assign img[11366] = 154;
assign img[11367] = 217;
assign img[11368] = 217;
assign img[11369] = 253;
assign img[11370] = 187;
assign img[11371] = 171;
assign img[11372] = 138;
assign img[11373] = 136;
assign img[11374] = 152;
assign img[11375] = 153;
assign img[11376] = 136;
assign img[11377] = 153;
assign img[11378] = 153;
assign img[11379] = 251;
assign img[11380] = 223;
assign img[11381] = 157;
assign img[11382] = 153;
assign img[11383] = 153;
assign img[11384] = 153;
assign img[11385] = 137;
assign img[11386] = 152;
assign img[11387] = 137;
assign img[11388] = 152;
assign img[11389] = 153;
assign img[11390] = 153;
assign img[11391] = 153;
assign img[11392] = 16;
assign img[11393] = 1;
assign img[11394] = 64;
assign img[11395] = 172;
assign img[11396] = 138;
assign img[11397] = 136;
assign img[11398] = 136;
assign img[11399] = 168;
assign img[11400] = 186;
assign img[11401] = 187;
assign img[11402] = 187;
assign img[11403] = 187;
assign img[11404] = 137;
assign img[11405] = 168;
assign img[11406] = 170;
assign img[11407] = 138;
assign img[11408] = 136;
assign img[11409] = 170;
assign img[11410] = 138;
assign img[11411] = 156;
assign img[11412] = 175;
assign img[11413] = 170;
assign img[11414] = 170;
assign img[11415] = 170;
assign img[11416] = 200;
assign img[11417] = 140;
assign img[11418] = 136;
assign img[11419] = 153;
assign img[11420] = 153;
assign img[11421] = 155;
assign img[11422] = 137;
assign img[11423] = 136;
assign img[11424] = 232;
assign img[11425] = 238;
assign img[11426] = 170;
assign img[11427] = 138;
assign img[11428] = 136;
assign img[11429] = 152;
assign img[11430] = 137;
assign img[11431] = 140;
assign img[11432] = 236;
assign img[11433] = 206;
assign img[11434] = 156;
assign img[11435] = 169;
assign img[11436] = 154;
assign img[11437] = 153;
assign img[11438] = 200;
assign img[11439] = 140;
assign img[11440] = 232;
assign img[11441] = 254;
assign img[11442] = 255;
assign img[11443] = 239;
assign img[11444] = 204;
assign img[11445] = 236;
assign img[11446] = 232;
assign img[11447] = 254;
assign img[11448] = 255;
assign img[11449] = 239;
assign img[11450] = 238;
assign img[11451] = 186;
assign img[11452] = 217;
assign img[11453] = 157;
assign img[11454] = 153;
assign img[11455] = 253;
assign img[11456] = 255;
assign img[11457] = 255;
assign img[11458] = 153;
assign img[11459] = 185;
assign img[11460] = 251;
assign img[11461] = 255;
assign img[11462] = 187;
assign img[11463] = 171;
assign img[11464] = 200;
assign img[11465] = 204;
assign img[11466] = 236;
assign img[11467] = 238;
assign img[11468] = 238;
assign img[11469] = 238;
assign img[11470] = 186;
assign img[11471] = 251;
assign img[11472] = 255;
assign img[11473] = 255;
assign img[11474] = 205;
assign img[11475] = 204;
assign img[11476] = 204;
assign img[11477] = 136;
assign img[11478] = 186;
assign img[11479] = 255;
assign img[11480] = 239;
assign img[11481] = 206;
assign img[11482] = 236;
assign img[11483] = 238;
assign img[11484] = 254;
assign img[11485] = 175;
assign img[11486] = 184;
assign img[11487] = 255;
assign img[11488] = 239;
assign img[11489] = 170;
assign img[11490] = 202;
assign img[11491] = 140;
assign img[11492] = 136;
assign img[11493] = 152;
assign img[11494] = 153;
assign img[11495] = 217;
assign img[11496] = 221;
assign img[11497] = 185;
assign img[11498] = 187;
assign img[11499] = 187;
assign img[11500] = 170;
assign img[11501] = 138;
assign img[11502] = 184;
assign img[11503] = 187;
assign img[11504] = 187;
assign img[11505] = 187;
assign img[11506] = 187;
assign img[11507] = 187;
assign img[11508] = 170;
assign img[11509] = 170;
assign img[11510] = 170;
assign img[11511] = 202;
assign img[11512] = 156;
assign img[11513] = 153;
assign img[11514] = 153;
assign img[11515] = 136;
assign img[11516] = 136;
assign img[11517] = 204;
assign img[11518] = 140;
assign img[11519] = 136;
assign img[11520] = 64;
assign img[11521] = 4;
assign img[11522] = 0;
assign img[11523] = 136;
assign img[11524] = 136;
assign img[11525] = 152;
assign img[11526] = 137;
assign img[11527] = 168;
assign img[11528] = 234;
assign img[11529] = 238;
assign img[11530] = 222;
assign img[11531] = 205;
assign img[11532] = 136;
assign img[11533] = 138;
assign img[11534] = 152;
assign img[11535] = 153;
assign img[11536] = 185;
assign img[11537] = 170;
assign img[11538] = 136;
assign img[11539] = 157;
assign img[11540] = 137;
assign img[11541] = 138;
assign img[11542] = 170;
assign img[11543] = 170;
assign img[11544] = 170;
assign img[11545] = 174;
assign img[11546] = 186;
assign img[11547] = 251;
assign img[11548] = 170;
assign img[11549] = 155;
assign img[11550] = 136;
assign img[11551] = 152;
assign img[11552] = 153;
assign img[11553] = 153;
assign img[11554] = 153;
assign img[11555] = 185;
assign img[11556] = 154;
assign img[11557] = 185;
assign img[11558] = 187;
assign img[11559] = 187;
assign img[11560] = 217;
assign img[11561] = 204;
assign img[11562] = 204;
assign img[11563] = 168;
assign img[11564] = 170;
assign img[11565] = 187;
assign img[11566] = 251;
assign img[11567] = 255;
assign img[11568] = 221;
assign img[11569] = 239;
assign img[11570] = 238;
assign img[11571] = 255;
assign img[11572] = 255;
assign img[11573] = 255;
assign img[11574] = 238;
assign img[11575] = 238;
assign img[11576] = 254;
assign img[11577] = 255;
assign img[11578] = 205;
assign img[11579] = 136;
assign img[11580] = 232;
assign img[11581] = 238;
assign img[11582] = 170;
assign img[11583] = 234;
assign img[11584] = 238;
assign img[11585] = 238;
assign img[11586] = 254;
assign img[11587] = 255;
assign img[11588] = 255;
assign img[11589] = 191;
assign img[11590] = 187;
assign img[11591] = 187;
assign img[11592] = 251;
assign img[11593] = 255;
assign img[11594] = 205;
assign img[11595] = 236;
assign img[11596] = 138;
assign img[11597] = 168;
assign img[11598] = 202;
assign img[11599] = 204;
assign img[11600] = 140;
assign img[11601] = 236;
assign img[11602] = 174;
assign img[11603] = 187;
assign img[11604] = 187;
assign img[11605] = 187;
assign img[11606] = 153;
assign img[11607] = 221;
assign img[11608] = 157;
assign img[11609] = 153;
assign img[11610] = 137;
assign img[11611] = 136;
assign img[11612] = 168;
assign img[11613] = 138;
assign img[11614] = 152;
assign img[11615] = 153;
assign img[11616] = 153;
assign img[11617] = 153;
assign img[11618] = 136;
assign img[11619] = 184;
assign img[11620] = 235;
assign img[11621] = 190;
assign img[11622] = 139;
assign img[11623] = 153;
assign img[11624] = 185;
assign img[11625] = 187;
assign img[11626] = 203;
assign img[11627] = 141;
assign img[11628] = 136;
assign img[11629] = 153;
assign img[11630] = 153;
assign img[11631] = 137;
assign img[11632] = 152;
assign img[11633] = 187;
assign img[11634] = 155;
assign img[11635] = 153;
assign img[11636] = 153;
assign img[11637] = 136;
assign img[11638] = 153;
assign img[11639] = 255;
assign img[11640] = 191;
assign img[11641] = 155;
assign img[11642] = 153;
assign img[11643] = 137;
assign img[11644] = 136;
assign img[11645] = 248;
assign img[11646] = 171;
assign img[11647] = 234;
assign img[11648] = 80;
assign img[11649] = 173;
assign img[11650] = 170;
assign img[11651] = 138;
assign img[11652] = 136;
assign img[11653] = 136;
assign img[11654] = 136;
assign img[11655] = 201;
assign img[11656] = 221;
assign img[11657] = 221;
assign img[11658] = 205;
assign img[11659] = 220;
assign img[11660] = 221;
assign img[11661] = 239;
assign img[11662] = 170;
assign img[11663] = 136;
assign img[11664] = 136;
assign img[11665] = 153;
assign img[11666] = 217;
assign img[11667] = 189;
assign img[11668] = 138;
assign img[11669] = 200;
assign img[11670] = 204;
assign img[11671] = 238;
assign img[11672] = 206;
assign img[11673] = 140;
assign img[11674] = 136;
assign img[11675] = 236;
assign img[11676] = 238;
assign img[11677] = 238;
assign img[11678] = 254;
assign img[11679] = 255;
assign img[11680] = 255;
assign img[11681] = 255;
assign img[11682] = 191;
assign img[11683] = 187;
assign img[11684] = 187;
assign img[11685] = 187;
assign img[11686] = 234;
assign img[11687] = 138;
assign img[11688] = 234;
assign img[11689] = 238;
assign img[11690] = 170;
assign img[11691] = 154;
assign img[11692] = 171;
assign img[11693] = 170;
assign img[11694] = 238;
assign img[11695] = 174;
assign img[11696] = 186;
assign img[11697] = 187;
assign img[11698] = 137;
assign img[11699] = 136;
assign img[11700] = 184;
assign img[11701] = 187;
assign img[11702] = 251;
assign img[11703] = 255;
assign img[11704] = 239;
assign img[11705] = 238;
assign img[11706] = 170;
assign img[11707] = 168;
assign img[11708] = 250;
assign img[11709] = 141;
assign img[11710] = 136;
assign img[11711] = 168;
assign img[11712] = 170;
assign img[11713] = 186;
assign img[11714] = 153;
assign img[11715] = 217;
assign img[11716] = 185;
assign img[11717] = 187;
assign img[11718] = 251;
assign img[11719] = 255;
assign img[11720] = 255;
assign img[11721] = 255;
assign img[11722] = 255;
assign img[11723] = 191;
assign img[11724] = 155;
assign img[11725] = 153;
assign img[11726] = 136;
assign img[11727] = 136;
assign img[11728] = 136;
assign img[11729] = 238;
assign img[11730] = 238;
assign img[11731] = 238;
assign img[11732] = 206;
assign img[11733] = 172;
assign img[11734] = 138;
assign img[11735] = 220;
assign img[11736] = 157;
assign img[11737] = 185;
assign img[11738] = 207;
assign img[11739] = 221;
assign img[11740] = 153;
assign img[11741] = 253;
assign img[11742] = 170;
assign img[11743] = 170;
assign img[11744] = 187;
assign img[11745] = 171;
assign img[11746] = 234;
assign img[11747] = 238;
assign img[11748] = 238;
assign img[11749] = 223;
assign img[11750] = 153;
assign img[11751] = 137;
assign img[11752] = 232;
assign img[11753] = 254;
assign img[11754] = 255;
assign img[11755] = 255;
assign img[11756] = 204;
assign img[11757] = 204;
assign img[11758] = 204;
assign img[11759] = 157;
assign img[11760] = 153;
assign img[11761] = 153;
assign img[11762] = 187;
assign img[11763] = 170;
assign img[11764] = 170;
assign img[11765] = 207;
assign img[11766] = 204;
assign img[11767] = 204;
assign img[11768] = 204;
assign img[11769] = 140;
assign img[11770] = 136;
assign img[11771] = 152;
assign img[11772] = 137;
assign img[11773] = 200;
assign img[11774] = 168;
assign img[11775] = 234;
assign img[11776] = 96;
assign img[11777] = 238;
assign img[11778] = 170;
assign img[11779] = 220;
assign img[11780] = 153;
assign img[11781] = 153;
assign img[11782] = 185;
assign img[11783] = 255;
assign img[11784] = 255;
assign img[11785] = 191;
assign img[11786] = 155;
assign img[11787] = 137;
assign img[11788] = 152;
assign img[11789] = 185;
assign img[11790] = 139;
assign img[11791] = 140;
assign img[11792] = 200;
assign img[11793] = 206;
assign img[11794] = 174;
assign img[11795] = 138;
assign img[11796] = 152;
assign img[11797] = 153;
assign img[11798] = 185;
assign img[11799] = 255;
assign img[11800] = 255;
assign img[11801] = 142;
assign img[11802] = 136;
assign img[11803] = 136;
assign img[11804] = 153;
assign img[11805] = 205;
assign img[11806] = 157;
assign img[11807] = 221;
assign img[11808] = 157;
assign img[11809] = 153;
assign img[11810] = 136;
assign img[11811] = 136;
assign img[11812] = 136;
assign img[11813] = 153;
assign img[11814] = 153;
assign img[11815] = 137;
assign img[11816] = 152;
assign img[11817] = 169;
assign img[11818] = 138;
assign img[11819] = 136;
assign img[11820] = 136;
assign img[11821] = 136;
assign img[11822] = 136;
assign img[11823] = 136;
assign img[11824] = 186;
assign img[11825] = 187;
assign img[11826] = 219;
assign img[11827] = 221;
assign img[11828] = 153;
assign img[11829] = 219;
assign img[11830] = 203;
assign img[11831] = 236;
assign img[11832] = 252;
assign img[11833] = 255;
assign img[11834] = 191;
assign img[11835] = 207;
assign img[11836] = 204;
assign img[11837] = 140;
assign img[11838] = 236;
assign img[11839] = 238;
assign img[11840] = 204;
assign img[11841] = 236;
assign img[11842] = 136;
assign img[11843] = 200;
assign img[11844] = 217;
assign img[11845] = 153;
assign img[11846] = 216;
assign img[11847] = 255;
assign img[11848] = 255;
assign img[11849] = 207;
assign img[11850] = 221;
assign img[11851] = 253;
assign img[11852] = 223;
assign img[11853] = 205;
assign img[11854] = 140;
assign img[11855] = 170;
assign img[11856] = 186;
assign img[11857] = 171;
assign img[11858] = 170;
assign img[11859] = 170;
assign img[11860] = 170;
assign img[11861] = 138;
assign img[11862] = 136;
assign img[11863] = 138;
assign img[11864] = 136;
assign img[11865] = 153;
assign img[11866] = 185;
assign img[11867] = 187;
assign img[11868] = 187;
assign img[11869] = 187;
assign img[11870] = 170;
assign img[11871] = 142;
assign img[11872] = 200;
assign img[11873] = 174;
assign img[11874] = 202;
assign img[11875] = 204;
assign img[11876] = 204;
assign img[11877] = 220;
assign img[11878] = 221;
assign img[11879] = 237;
assign img[11880] = 238;
assign img[11881] = 174;
assign img[11882] = 184;
assign img[11883] = 159;
assign img[11884] = 137;
assign img[11885] = 168;
assign img[11886] = 234;
assign img[11887] = 254;
assign img[11888] = 223;
assign img[11889] = 221;
assign img[11890] = 136;
assign img[11891] = 153;
assign img[11892] = 153;
assign img[11893] = 153;
assign img[11894] = 153;
assign img[11895] = 251;
assign img[11896] = 255;
assign img[11897] = 255;
assign img[11898] = 127;
assign img[11899] = 7;
assign img[11900] = 34;
assign img[11901] = 226;
assign img[11902] = 238;
assign img[11903] = 238;
assign img[11904] = 96;
assign img[11905] = 238;
assign img[11906] = 238;
assign img[11907] = 206;
assign img[11908] = 204;
assign img[11909] = 140;
assign img[11910] = 168;
assign img[11911] = 191;
assign img[11912] = 187;
assign img[11913] = 175;
assign img[11914] = 170;
assign img[11915] = 170;
assign img[11916] = 152;
assign img[11917] = 153;
assign img[11918] = 187;
assign img[11919] = 171;
assign img[11920] = 186;
assign img[11921] = 191;
assign img[11922] = 255;
assign img[11923] = 255;
assign img[11924] = 255;
assign img[11925] = 187;
assign img[11926] = 187;
assign img[11927] = 187;
assign img[11928] = 234;
assign img[11929] = 174;
assign img[11930] = 136;
assign img[11931] = 136;
assign img[11932] = 204;
assign img[11933] = 236;
assign img[11934] = 254;
assign img[11935] = 159;
assign img[11936] = 153;
assign img[11937] = 153;
assign img[11938] = 153;
assign img[11939] = 153;
assign img[11940] = 153;
assign img[11941] = 136;
assign img[11942] = 200;
assign img[11943] = 156;
assign img[11944] = 187;
assign img[11945] = 155;
assign img[11946] = 136;
assign img[11947] = 152;
assign img[11948] = 153;
assign img[11949] = 153;
assign img[11950] = 232;
assign img[11951] = 255;
assign img[11952] = 255;
assign img[11953] = 255;
assign img[11954] = 255;
assign img[11955] = 175;
assign img[11956] = 170;
assign img[11957] = 238;
assign img[11958] = 254;
assign img[11959] = 255;
assign img[11960] = 255;
assign img[11961] = 255;
assign img[11962] = 155;
assign img[11963] = 153;
assign img[11964] = 185;
assign img[11965] = 155;
assign img[11966] = 137;
assign img[11967] = 153;
assign img[11968] = 153;
assign img[11969] = 153;
assign img[11970] = 200;
assign img[11971] = 168;
assign img[11972] = 170;
assign img[11973] = 154;
assign img[11974] = 136;
assign img[11975] = 153;
assign img[11976] = 200;
assign img[11977] = 236;
assign img[11978] = 206;
assign img[11979] = 204;
assign img[11980] = 136;
assign img[11981] = 250;
assign img[11982] = 255;
assign img[11983] = 223;
assign img[11984] = 204;
assign img[11985] = 238;
assign img[11986] = 174;
assign img[11987] = 186;
assign img[11988] = 153;
assign img[11989] = 153;
assign img[11990] = 136;
assign img[11991] = 168;
assign img[11992] = 170;
assign img[11993] = 234;
assign img[11994] = 220;
assign img[11995] = 140;
assign img[11996] = 184;
assign img[11997] = 155;
assign img[11998] = 185;
assign img[11999] = 223;
assign img[12000] = 136;
assign img[12001] = 168;
assign img[12002] = 234;
assign img[12003] = 239;
assign img[12004] = 255;
assign img[12005] = 223;
assign img[12006] = 185;
assign img[12007] = 251;
assign img[12008] = 187;
assign img[12009] = 255;
assign img[12010] = 187;
assign img[12011] = 187;
assign img[12012] = 187;
assign img[12013] = 251;
assign img[12014] = 255;
assign img[12015] = 239;
assign img[12016] = 140;
assign img[12017] = 136;
assign img[12018] = 168;
assign img[12019] = 170;
assign img[12020] = 170;
assign img[12021] = 170;
assign img[12022] = 170;
assign img[12023] = 186;
assign img[12024] = 251;
assign img[12025] = 255;
assign img[12026] = 187;
assign img[12027] = 187;
assign img[12028] = 137;
assign img[12029] = 232;
assign img[12030] = 238;
assign img[12031] = 255;
assign img[12032] = 96;
assign img[12033] = 238;
assign img[12034] = 238;
assign img[12035] = 206;
assign img[12036] = 152;
assign img[12037] = 187;
assign img[12038] = 187;
assign img[12039] = 171;
assign img[12040] = 234;
assign img[12041] = 239;
assign img[12042] = 238;
assign img[12043] = 170;
assign img[12044] = 170;
assign img[12045] = 170;
assign img[12046] = 170;
assign img[12047] = 170;
assign img[12048] = 170;
assign img[12049] = 170;
assign img[12050] = 250;
assign img[12051] = 255;
assign img[12052] = 170;
assign img[12053] = 170;
assign img[12054] = 170;
assign img[12055] = 187;
assign img[12056] = 153;
assign img[12057] = 153;
assign img[12058] = 169;
assign img[12059] = 238;
assign img[12060] = 206;
assign img[12061] = 238;
assign img[12062] = 174;
assign img[12063] = 170;
assign img[12064] = 136;
assign img[12065] = 236;
assign img[12066] = 238;
assign img[12067] = 238;
assign img[12068] = 204;
assign img[12069] = 221;
assign img[12070] = 221;
assign img[12071] = 221;
assign img[12072] = 153;
assign img[12073] = 201;
assign img[12074] = 168;
assign img[12075] = 170;
assign img[12076] = 170;
assign img[12077] = 138;
assign img[12078] = 136;
assign img[12079] = 136;
assign img[12080] = 232;
assign img[12081] = 239;
assign img[12082] = 238;
assign img[12083] = 238;
assign img[12084] = 186;
assign img[12085] = 251;
assign img[12086] = 187;
assign img[12087] = 187;
assign img[12088] = 171;
assign img[12089] = 206;
assign img[12090] = 204;
assign img[12091] = 205;
assign img[12092] = 204;
assign img[12093] = 136;
assign img[12094] = 152;
assign img[12095] = 233;
assign img[12096] = 238;
assign img[12097] = 238;
assign img[12098] = 204;
assign img[12099] = 252;
assign img[12100] = 239;
assign img[12101] = 190;
assign img[12102] = 238;
assign img[12103] = 238;
assign img[12104] = 136;
assign img[12105] = 152;
assign img[12106] = 249;
assign img[12107] = 190;
assign img[12108] = 187;
assign img[12109] = 187;
assign img[12110] = 235;
assign img[12111] = 238;
assign img[12112] = 254;
assign img[12113] = 255;
assign img[12114] = 223;
assign img[12115] = 157;
assign img[12116] = 153;
assign img[12117] = 187;
assign img[12118] = 187;
assign img[12119] = 187;
assign img[12120] = 187;
assign img[12121] = 255;
assign img[12122] = 238;
assign img[12123] = 223;
assign img[12124] = 221;
assign img[12125] = 253;
assign img[12126] = 238;
assign img[12127] = 207;
assign img[12128] = 220;
assign img[12129] = 189;
assign img[12130] = 251;
assign img[12131] = 207;
assign img[12132] = 220;
assign img[12133] = 221;
assign img[12134] = 136;
assign img[12135] = 184;
assign img[12136] = 202;
assign img[12137] = 253;
assign img[12138] = 187;
assign img[12139] = 187;
assign img[12140] = 169;
assign img[12141] = 234;
assign img[12142] = 254;
assign img[12143] = 239;
assign img[12144] = 238;
assign img[12145] = 238;
assign img[12146] = 238;
assign img[12147] = 170;
assign img[12148] = 186;
assign img[12149] = 155;
assign img[12150] = 168;
assign img[12151] = 238;
assign img[12152] = 238;
assign img[12153] = 238;
assign img[12154] = 174;
assign img[12155] = 170;
assign img[12156] = 152;
assign img[12157] = 249;
assign img[12158] = 255;
assign img[12159] = 255;
assign img[12160] = 64;
assign img[12161] = 68;
assign img[12162] = 68;
assign img[12163] = 254;
assign img[12164] = 239;
assign img[12165] = 174;
assign img[12166] = 204;
assign img[12167] = 236;
assign img[12168] = 238;
assign img[12169] = 239;
assign img[12170] = 238;
assign img[12171] = 238;
assign img[12172] = 238;
assign img[12173] = 174;
assign img[12174] = 186;
assign img[12175] = 187;
assign img[12176] = 187;
assign img[12177] = 239;
assign img[12178] = 238;
assign img[12179] = 174;
assign img[12180] = 170;
assign img[12181] = 187;
assign img[12182] = 171;
assign img[12183] = 202;
assign img[12184] = 238;
assign img[12185] = 159;
assign img[12186] = 153;
assign img[12187] = 155;
assign img[12188] = 185;
assign img[12189] = 255;
assign img[12190] = 204;
assign img[12191] = 238;
assign img[12192] = 76;
assign img[12193] = 228;
assign img[12194] = 191;
assign img[12195] = 255;
assign img[12196] = 157;
assign img[12197] = 153;
assign img[12198] = 153;
assign img[12199] = 153;
assign img[12200] = 201;
assign img[12201] = 221;
assign img[12202] = 137;
assign img[12203] = 170;
assign img[12204] = 170;
assign img[12205] = 170;
assign img[12206] = 250;
assign img[12207] = 191;
assign img[12208] = 187;
assign img[12209] = 187;
assign img[12210] = 155;
assign img[12211] = 157;
assign img[12212] = 221;
assign img[12213] = 223;
assign img[12214] = 205;
assign img[12215] = 204;
assign img[12216] = 252;
assign img[12217] = 255;
assign img[12218] = 207;
assign img[12219] = 188;
assign img[12220] = 251;
assign img[12221] = 191;
assign img[12222] = 155;
assign img[12223] = 153;
assign img[12224] = 153;
assign img[12225] = 139;
assign img[12226] = 170;
assign img[12227] = 234;
assign img[12228] = 174;
assign img[12229] = 138;
assign img[12230] = 152;
assign img[12231] = 191;
assign img[12232] = 255;
assign img[12233] = 255;
assign img[12234] = 255;
assign img[12235] = 239;
assign img[12236] = 254;
assign img[12237] = 207;
assign img[12238] = 236;
assign img[12239] = 255;
assign img[12240] = 238;
assign img[12241] = 238;
assign img[12242] = 238;
assign img[12243] = 255;
assign img[12244] = 255;
assign img[12245] = 255;
assign img[12246] = 238;
assign img[12247] = 239;
assign img[12248] = 191;
assign img[12249] = 171;
assign img[12250] = 152;
assign img[12251] = 185;
assign img[12252] = 170;
assign img[12253] = 168;
assign img[12254] = 234;
assign img[12255] = 238;
assign img[12256] = 136;
assign img[12257] = 157;
assign img[12258] = 239;
assign img[12259] = 223;
assign img[12260] = 221;
assign img[12261] = 221;
assign img[12262] = 153;
assign img[12263] = 249;
assign img[12264] = 223;
assign img[12265] = 253;
assign img[12266] = 238;
assign img[12267] = 174;
assign img[12268] = 170;
assign img[12269] = 234;
assign img[12270] = 238;
assign img[12271] = 254;
assign img[12272] = 157;
assign img[12273] = 153;
assign img[12274] = 217;
assign img[12275] = 221;
assign img[12276] = 253;
assign img[12277] = 255;
assign img[12278] = 239;
assign img[12279] = 238;
assign img[12280] = 238;
assign img[12281] = 222;
assign img[12282] = 253;
assign img[12283] = 191;
assign img[12284] = 170;
assign img[12285] = 238;
assign img[12286] = 238;
assign img[12287] = 254;
assign img[12288] = 96;
assign img[12289] = 238;
assign img[12290] = 238;
assign img[12291] = 255;
assign img[12292] = 255;
assign img[12293] = 191;
assign img[12294] = 187;
assign img[12295] = 187;
assign img[12296] = 251;
assign img[12297] = 223;
assign img[12298] = 221;
assign img[12299] = 255;
assign img[12300] = 155;
assign img[12301] = 153;
assign img[12302] = 217;
assign img[12303] = 189;
assign img[12304] = 251;
assign img[12305] = 191;
assign img[12306] = 221;
assign img[12307] = 253;
assign img[12308] = 171;
assign img[12309] = 170;
assign img[12310] = 186;
assign img[12311] = 255;
assign img[12312] = 191;
assign img[12313] = 187;
assign img[12314] = 170;
assign img[12315] = 170;
assign img[12316] = 170;
assign img[12317] = 238;
assign img[12318] = 238;
assign img[12319] = 238;
assign img[12320] = 152;
assign img[12321] = 249;
assign img[12322] = 223;
assign img[12323] = 205;
assign img[12324] = 204;
assign img[12325] = 168;
assign img[12326] = 170;
assign img[12327] = 170;
assign img[12328] = 170;
assign img[12329] = 255;
assign img[12330] = 191;
assign img[12331] = 187;
assign img[12332] = 171;
assign img[12333] = 170;
assign img[12334] = 234;
assign img[12335] = 174;
assign img[12336] = 186;
assign img[12337] = 139;
assign img[12338] = 136;
assign img[12339] = 251;
assign img[12340] = 187;
assign img[12341] = 187;
assign img[12342] = 251;
assign img[12343] = 239;
assign img[12344] = 170;
assign img[12345] = 251;
assign img[12346] = 137;
assign img[12347] = 152;
assign img[12348] = 169;
assign img[12349] = 174;
assign img[12350] = 238;
assign img[12351] = 138;
assign img[12352] = 216;
assign img[12353] = 253;
assign img[12354] = 255;
assign img[12355] = 187;
assign img[12356] = 170;
assign img[12357] = 171;
assign img[12358] = 234;
assign img[12359] = 191;
assign img[12360] = 171;
assign img[12361] = 234;
assign img[12362] = 170;
assign img[12363] = 170;
assign img[12364] = 170;
assign img[12365] = 187;
assign img[12366] = 251;
assign img[12367] = 255;
assign img[12368] = 191;
assign img[12369] = 251;
assign img[12370] = 191;
assign img[12371] = 187;
assign img[12372] = 187;
assign img[12373] = 187;
assign img[12374] = 234;
assign img[12375] = 238;
assign img[12376] = 238;
assign img[12377] = 170;
assign img[12378] = 170;
assign img[12379] = 186;
assign img[12380] = 153;
assign img[12381] = 157;
assign img[12382] = 253;
assign img[12383] = 191;
assign img[12384] = 187;
assign img[12385] = 187;
assign img[12386] = 251;
assign img[12387] = 239;
assign img[12388] = 238;
assign img[12389] = 238;
assign img[12390] = 170;
assign img[12391] = 170;
assign img[12392] = 234;
assign img[12393] = 238;
assign img[12394] = 186;
assign img[12395] = 187;
assign img[12396] = 170;
assign img[12397] = 202;
assign img[12398] = 184;
assign img[12399] = 187;
assign img[12400] = 187;
assign img[12401] = 170;
assign img[12402] = 138;
assign img[12403] = 136;
assign img[12404] = 184;
assign img[12405] = 187;
assign img[12406] = 187;
assign img[12407] = 255;
assign img[12408] = 191;
assign img[12409] = 155;
assign img[12410] = 153;
assign img[12411] = 187;
assign img[12412] = 187;
assign img[12413] = 251;
assign img[12414] = 255;
assign img[12415] = 255;
assign img[12416] = 64;
assign img[12417] = 204;
assign img[12418] = 236;
assign img[12419] = 255;
assign img[12420] = 206;
assign img[12421] = 204;
assign img[12422] = 204;
assign img[12423] = 204;
assign img[12424] = 220;
assign img[12425] = 221;
assign img[12426] = 221;
assign img[12427] = 253;
assign img[12428] = 255;
assign img[12429] = 223;
assign img[12430] = 137;
assign img[12431] = 136;
assign img[12432] = 216;
assign img[12433] = 221;
assign img[12434] = 205;
assign img[12435] = 220;
assign img[12436] = 185;
assign img[12437] = 251;
assign img[12438] = 223;
assign img[12439] = 221;
assign img[12440] = 140;
assign img[12441] = 137;
assign img[12442] = 136;
assign img[12443] = 136;
assign img[12444] = 200;
assign img[12445] = 204;
assign img[12446] = 204;
assign img[12447] = 236;
assign img[12448] = 206;
assign img[12449] = 236;
assign img[12450] = 238;
assign img[12451] = 238;
assign img[12452] = 142;
assign img[12453] = 153;
assign img[12454] = 201;
assign img[12455] = 204;
assign img[12456] = 204;
assign img[12457] = 204;
assign img[12458] = 254;
assign img[12459] = 155;
assign img[12460] = 153;
assign img[12461] = 139;
assign img[12462] = 232;
assign img[12463] = 238;
assign img[12464] = 238;
assign img[12465] = 255;
assign img[12466] = 251;
assign img[12467] = 191;
assign img[12468] = 255;
assign img[12469] = 191;
assign img[12470] = 187;
assign img[12471] = 223;
assign img[12472] = 253;
assign img[12473] = 221;
assign img[12474] = 157;
assign img[12475] = 153;
assign img[12476] = 153;
assign img[12477] = 153;
assign img[12478] = 153;
assign img[12479] = 137;
assign img[12480] = 216;
assign img[12481] = 157;
assign img[12482] = 185;
assign img[12483] = 139;
assign img[12484] = 170;
assign img[12485] = 171;
assign img[12486] = 170;
assign img[12487] = 170;
assign img[12488] = 216;
assign img[12489] = 221;
assign img[12490] = 253;
assign img[12491] = 255;
assign img[12492] = 255;
assign img[12493] = 191;
assign img[12494] = 187;
assign img[12495] = 251;
assign img[12496] = 187;
assign img[12497] = 251;
assign img[12498] = 255;
assign img[12499] = 187;
assign img[12500] = 155;
assign img[12501] = 153;
assign img[12502] = 234;
assign img[12503] = 204;
assign img[12504] = 204;
assign img[12505] = 204;
assign img[12506] = 140;
assign img[12507] = 157;
assign img[12508] = 185;
assign img[12509] = 187;
assign img[12510] = 251;
assign img[12511] = 223;
assign img[12512] = 253;
assign img[12513] = 255;
assign img[12514] = 238;
assign img[12515] = 206;
assign img[12516] = 220;
assign img[12517] = 157;
assign img[12518] = 153;
assign img[12519] = 153;
assign img[12520] = 217;
assign img[12521] = 205;
assign img[12522] = 236;
assign img[12523] = 174;
assign img[12524] = 138;
assign img[12525] = 200;
assign img[12526] = 204;
assign img[12527] = 206;
assign img[12528] = 174;
assign img[12529] = 170;
assign img[12530] = 154;
assign img[12531] = 185;
assign img[12532] = 187;
assign img[12533] = 235;
assign img[12534] = 254;
assign img[12535] = 255;
assign img[12536] = 223;
assign img[12537] = 221;
assign img[12538] = 221;
assign img[12539] = 159;
assign img[12540] = 171;
assign img[12541] = 238;
assign img[12542] = 254;
assign img[12543] = 255;
assign img[12544] = 96;
assign img[12545] = 239;
assign img[12546] = 238;
assign img[12547] = 191;
assign img[12548] = 171;
assign img[12549] = 186;
assign img[12550] = 251;
assign img[12551] = 255;
assign img[12552] = 255;
assign img[12553] = 255;
assign img[12554] = 223;
assign img[12555] = 255;
assign img[12556] = 187;
assign img[12557] = 187;
assign img[12558] = 153;
assign img[12559] = 153;
assign img[12560] = 137;
assign img[12561] = 136;
assign img[12562] = 184;
assign img[12563] = 251;
assign img[12564] = 255;
assign img[12565] = 255;
assign img[12566] = 239;
assign img[12567] = 255;
assign img[12568] = 255;
assign img[12569] = 191;
assign img[12570] = 153;
assign img[12571] = 205;
assign img[12572] = 236;
assign img[12573] = 238;
assign img[12574] = 190;
assign img[12575] = 187;
assign img[12576] = 187;
assign img[12577] = 187;
assign img[12578] = 138;
assign img[12579] = 238;
assign img[12580] = 174;
assign img[12581] = 170;
assign img[12582] = 170;
assign img[12583] = 155;
assign img[12584] = 217;
assign img[12585] = 221;
assign img[12586] = 221;
assign img[12587] = 191;
assign img[12588] = 187;
assign img[12589] = 187;
assign img[12590] = 255;
assign img[12591] = 239;
assign img[12592] = 154;
assign img[12593] = 205;
assign img[12594] = 204;
assign img[12595] = 172;
assign img[12596] = 234;
assign img[12597] = 255;
assign img[12598] = 191;
assign img[12599] = 187;
assign img[12600] = 153;
assign img[12601] = 187;
assign img[12602] = 187;
assign img[12603] = 139;
assign img[12604] = 136;
assign img[12605] = 153;
assign img[12606] = 201;
assign img[12607] = 236;
assign img[12608] = 238;
assign img[12609] = 206;
assign img[12610] = 140;
assign img[12611] = 255;
assign img[12612] = 223;
assign img[12613] = 157;
assign img[12614] = 153;
assign img[12615] = 153;
assign img[12616] = 153;
assign img[12617] = 187;
assign img[12618] = 219;
assign img[12619] = 221;
assign img[12620] = 153;
assign img[12621] = 219;
assign img[12622] = 187;
assign img[12623] = 223;
assign img[12624] = 253;
assign img[12625] = 255;
assign img[12626] = 255;
assign img[12627] = 255;
assign img[12628] = 238;
assign img[12629] = 238;
assign img[12630] = 136;
assign img[12631] = 204;
assign img[12632] = 238;
assign img[12633] = 191;
assign img[12634] = 187;
assign img[12635] = 187;
assign img[12636] = 234;
assign img[12637] = 255;
assign img[12638] = 171;
assign img[12639] = 174;
assign img[12640] = 170;
assign img[12641] = 170;
assign img[12642] = 250;
assign img[12643] = 255;
assign img[12644] = 187;
assign img[12645] = 191;
assign img[12646] = 139;
assign img[12647] = 204;
assign img[12648] = 236;
assign img[12649] = 239;
assign img[12650] = 238;
assign img[12651] = 238;
assign img[12652] = 170;
assign img[12653] = 170;
assign img[12654] = 251;
assign img[12655] = 239;
assign img[12656] = 255;
assign img[12657] = 153;
assign img[12658] = 153;
assign img[12659] = 185;
assign img[12660] = 187;
assign img[12661] = 187;
assign img[12662] = 187;
assign img[12663] = 255;
assign img[12664] = 255;
assign img[12665] = 159;
assign img[12666] = 153;
assign img[12667] = 137;
assign img[12668] = 168;
assign img[12669] = 234;
assign img[12670] = 206;
assign img[12671] = 238;
assign img[12672] = 96;
assign img[12673] = 255;
assign img[12674] = 255;
assign img[12675] = 191;
assign img[12676] = 155;
assign img[12677] = 187;
assign img[12678] = 155;
assign img[12679] = 136;
assign img[12680] = 200;
assign img[12681] = 220;
assign img[12682] = 221;
assign img[12683] = 237;
assign img[12684] = 238;
assign img[12685] = 236;
assign img[12686] = 136;
assign img[12687] = 170;
assign img[12688] = 136;
assign img[12689] = 136;
assign img[12690] = 200;
assign img[12691] = 142;
assign img[12692] = 136;
assign img[12693] = 238;
assign img[12694] = 158;
assign img[12695] = 201;
assign img[12696] = 204;
assign img[12697] = 140;
assign img[12698] = 136;
assign img[12699] = 204;
assign img[12700] = 204;
assign img[12701] = 206;
assign img[12702] = 238;
assign img[12703] = 238;
assign img[12704] = 238;
assign img[12705] = 238;
assign img[12706] = 238;
assign img[12707] = 170;
assign img[12708] = 186;
assign img[12709] = 153;
assign img[12710] = 185;
assign img[12711] = 187;
assign img[12712] = 219;
assign img[12713] = 205;
assign img[12714] = 136;
assign img[12715] = 185;
assign img[12716] = 187;
assign img[12717] = 171;
assign img[12718] = 250;
assign img[12719] = 239;
assign img[12720] = 170;
assign img[12721] = 171;
assign img[12722] = 170;
assign img[12723] = 170;
assign img[12724] = 170;
assign img[12725] = 234;
assign img[12726] = 238;
assign img[12727] = 170;
assign img[12728] = 170;
assign img[12729] = 170;
assign img[12730] = 136;
assign img[12731] = 137;
assign img[12732] = 234;
assign img[12733] = 206;
assign img[12734] = 236;
assign img[12735] = 239;
assign img[12736] = 238;
assign img[12737] = 254;
assign img[12738] = 239;
assign img[12739] = 238;
assign img[12740] = 238;
assign img[12741] = 190;
assign img[12742] = 187;
assign img[12743] = 191;
assign img[12744] = 170;
assign img[12745] = 170;
assign img[12746] = 186;
assign img[12747] = 187;
assign img[12748] = 187;
assign img[12749] = 171;
assign img[12750] = 170;
assign img[12751] = 186;
assign img[12752] = 187;
assign img[12753] = 223;
assign img[12754] = 221;
assign img[12755] = 153;
assign img[12756] = 185;
assign img[12757] = 155;
assign img[12758] = 137;
assign img[12759] = 204;
assign img[12760] = 140;
assign img[12761] = 174;
assign img[12762] = 138;
assign img[12763] = 136;
assign img[12764] = 185;
assign img[12765] = 171;
assign img[12766] = 234;
assign img[12767] = 174;
assign img[12768] = 186;
assign img[12769] = 187;
assign img[12770] = 251;
assign img[12771] = 255;
assign img[12772] = 155;
assign img[12773] = 153;
assign img[12774] = 155;
assign img[12775] = 171;
assign img[12776] = 186;
assign img[12777] = 187;
assign img[12778] = 250;
assign img[12779] = 255;
assign img[12780] = 155;
assign img[12781] = 217;
assign img[12782] = 153;
assign img[12783] = 153;
assign img[12784] = 153;
assign img[12785] = 185;
assign img[12786] = 187;
assign img[12787] = 185;
assign img[12788] = 187;
assign img[12789] = 187;
assign img[12790] = 217;
assign img[12791] = 239;
assign img[12792] = 206;
assign img[12793] = 206;
assign img[12794] = 204;
assign img[12795] = 142;
assign img[12796] = 168;
assign img[12797] = 234;
assign img[12798] = 238;
assign img[12799] = 238;
assign img[12800] = 96;
assign img[12801] = 239;
assign img[12802] = 238;
assign img[12803] = 223;
assign img[12804] = 204;
assign img[12805] = 204;
assign img[12806] = 220;
assign img[12807] = 205;
assign img[12808] = 236;
assign img[12809] = 238;
assign img[12810] = 204;
assign img[12811] = 238;
assign img[12812] = 186;
assign img[12813] = 255;
assign img[12814] = 157;
assign img[12815] = 153;
assign img[12816] = 201;
assign img[12817] = 204;
assign img[12818] = 204;
assign img[12819] = 238;
assign img[12820] = 238;
assign img[12821] = 238;
assign img[12822] = 254;
assign img[12823] = 239;
assign img[12824] = 238;
assign img[12825] = 238;
assign img[12826] = 238;
assign img[12827] = 238;
assign img[12828] = 238;
assign img[12829] = 254;
assign img[12830] = 255;
assign img[12831] = 191;
assign img[12832] = 136;
assign img[12833] = 254;
assign img[12834] = 207;
assign img[12835] = 204;
assign img[12836] = 221;
assign img[12837] = 221;
assign img[12838] = 204;
assign img[12839] = 204;
assign img[12840] = 204;
assign img[12841] = 204;
assign img[12842] = 204;
assign img[12843] = 238;
assign img[12844] = 254;
assign img[12845] = 175;
assign img[12846] = 234;
assign img[12847] = 238;
assign img[12848] = 238;
assign img[12849] = 206;
assign img[12850] = 204;
assign img[12851] = 204;
assign img[12852] = 184;
assign img[12853] = 251;
assign img[12854] = 255;
assign img[12855] = 238;
assign img[12856] = 170;
assign img[12857] = 171;
assign img[12858] = 187;
assign img[12859] = 251;
assign img[12860] = 221;
assign img[12861] = 157;
assign img[12862] = 153;
assign img[12863] = 249;
assign img[12864] = 255;
assign img[12865] = 191;
assign img[12866] = 187;
assign img[12867] = 187;
assign img[12868] = 251;
assign img[12869] = 191;
assign img[12870] = 187;
assign img[12871] = 187;
assign img[12872] = 187;
assign img[12873] = 187;
assign img[12874] = 251;
assign img[12875] = 191;
assign img[12876] = 171;
assign img[12877] = 170;
assign img[12878] = 186;
assign img[12879] = 255;
assign img[12880] = 255;
assign img[12881] = 239;
assign img[12882] = 174;
assign img[12883] = 170;
assign img[12884] = 234;
assign img[12885] = 238;
assign img[12886] = 220;
assign img[12887] = 221;
assign img[12888] = 204;
assign img[12889] = 204;
assign img[12890] = 204;
assign img[12891] = 204;
assign img[12892] = 152;
assign img[12893] = 205;
assign img[12894] = 252;
assign img[12895] = 255;
assign img[12896] = 155;
assign img[12897] = 185;
assign img[12898] = 187;
assign img[12899] = 171;
assign img[12900] = 234;
assign img[12901] = 223;
assign img[12902] = 153;
assign img[12903] = 187;
assign img[12904] = 187;
assign img[12905] = 191;
assign img[12906] = 255;
assign img[12907] = 239;
assign img[12908] = 238;
assign img[12909] = 238;
assign img[12910] = 254;
assign img[12911] = 255;
assign img[12912] = 157;
assign img[12913] = 185;
assign img[12914] = 251;
assign img[12915] = 255;
assign img[12916] = 239;
assign img[12917] = 238;
assign img[12918] = 238;
assign img[12919] = 238;
assign img[12920] = 238;
assign img[12921] = 238;
assign img[12922] = 221;
assign img[12923] = 205;
assign img[12924] = 204;
assign img[12925] = 236;
assign img[12926] = 238;
assign img[12927] = 238;
assign img[12928] = 0;
assign img[12929] = 230;
assign img[12930] = 206;
assign img[12931] = 204;
assign img[12932] = 236;
assign img[12933] = 191;
assign img[12934] = 175;
assign img[12935] = 138;
assign img[12936] = 238;
assign img[12937] = 206;
assign img[12938] = 238;
assign img[12939] = 239;
assign img[12940] = 206;
assign img[12941] = 204;
assign img[12942] = 252;
assign img[12943] = 187;
assign img[12944] = 187;
assign img[12945] = 187;
assign img[12946] = 187;
assign img[12947] = 187;
assign img[12948] = 187;
assign img[12949] = 251;
assign img[12950] = 187;
assign img[12951] = 187;
assign img[12952] = 187;
assign img[12953] = 187;
assign img[12954] = 187;
assign img[12955] = 217;
assign img[12956] = 204;
assign img[12957] = 204;
assign img[12958] = 252;
assign img[12959] = 191;
assign img[12960] = 136;
assign img[12961] = 136;
assign img[12962] = 168;
assign img[12963] = 251;
assign img[12964] = 171;
assign img[12965] = 170;
assign img[12966] = 234;
assign img[12967] = 238;
assign img[12968] = 110;
assign img[12969] = 86;
assign img[12970] = 100;
assign img[12971] = 149;
assign img[12972] = 153;
assign img[12973] = 153;
assign img[12974] = 232;
assign img[12975] = 238;
assign img[12976] = 238;
assign img[12977] = 239;
assign img[12978] = 255;
assign img[12979] = 170;
assign img[12980] = 170;
assign img[12981] = 234;
assign img[12982] = 204;
assign img[12983] = 204;
assign img[12984] = 204;
assign img[12985] = 204;
assign img[12986] = 204;
assign img[12987] = 204;
assign img[12988] = 221;
assign img[12989] = 157;
assign img[12990] = 137;
assign img[12991] = 234;
assign img[12992] = 238;
assign img[12993] = 175;
assign img[12994] = 170;
assign img[12995] = 234;
assign img[12996] = 202;
assign img[12997] = 204;
assign img[12998] = 220;
assign img[12999] = 221;
assign img[13000] = 205;
assign img[13001] = 204;
assign img[13002] = 220;
assign img[13003] = 237;
assign img[13004] = 138;
assign img[13005] = 170;
assign img[13006] = 250;
assign img[13007] = 255;
assign img[13008] = 255;
assign img[13009] = 255;
assign img[13010] = 174;
assign img[13011] = 174;
assign img[13012] = 154;
assign img[13013] = 155;
assign img[13014] = 153;
assign img[13015] = 221;
assign img[13016] = 253;
assign img[13017] = 223;
assign img[13018] = 157;
assign img[13019] = 187;
assign img[13020] = 138;
assign img[13021] = 153;
assign img[13022] = 153;
assign img[13023] = 153;
assign img[13024] = 153;
assign img[13025] = 185;
assign img[13026] = 251;
assign img[13027] = 223;
assign img[13028] = 204;
assign img[13029] = 220;
assign img[13030] = 221;
assign img[13031] = 185;
assign img[13032] = 171;
assign img[13033] = 187;
assign img[13034] = 251;
assign img[13035] = 191;
assign img[13036] = 138;
assign img[13037] = 251;
assign img[13038] = 139;
assign img[13039] = 168;
assign img[13040] = 170;
assign img[13041] = 170;
assign img[13042] = 170;
assign img[13043] = 202;
assign img[13044] = 172;
assign img[13045] = 218;
assign img[13046] = 221;
assign img[13047] = 255;
assign img[13048] = 255;
assign img[13049] = 239;
assign img[13050] = 238;
assign img[13051] = 174;
assign img[13052] = 202;
assign img[13053] = 204;
assign img[13054] = 236;
assign img[13055] = 239;
assign img[13056] = 96;
assign img[13057] = 191;
assign img[13058] = 235;
assign img[13059] = 239;
assign img[13060] = 168;
assign img[13061] = 139;
assign img[13062] = 136;
assign img[13063] = 201;
assign img[13064] = 236;
assign img[13065] = 238;
assign img[13066] = 254;
assign img[13067] = 255;
assign img[13068] = 239;
assign img[13069] = 238;
assign img[13070] = 238;
assign img[13071] = 255;
assign img[13072] = 255;
assign img[13073] = 191;
assign img[13074] = 219;
assign img[13075] = 157;
assign img[13076] = 153;
assign img[13077] = 217;
assign img[13078] = 201;
assign img[13079] = 236;
assign img[13080] = 255;
assign img[13081] = 175;
assign img[13082] = 254;
assign img[13083] = 255;
assign img[13084] = 255;
assign img[13085] = 255;
assign img[13086] = 191;
assign img[13087] = 171;
assign img[13088] = 136;
assign img[13089] = 136;
assign img[13090] = 136;
assign img[13091] = 234;
assign img[13092] = 204;
assign img[13093] = 236;
assign img[13094] = 170;
assign img[13095] = 187;
assign img[13096] = 234;
assign img[13097] = 206;
assign img[13098] = 136;
assign img[13099] = 170;
assign img[13100] = 186;
assign img[13101] = 239;
assign img[13102] = 238;
assign img[13103] = 238;
assign img[13104] = 238;
assign img[13105] = 191;
assign img[13106] = 255;
assign img[13107] = 187;
assign img[13108] = 170;
assign img[13109] = 250;
assign img[13110] = 255;
assign img[13111] = 206;
assign img[13112] = 204;
assign img[13113] = 172;
assign img[13114] = 170;
assign img[13115] = 157;
assign img[13116] = 255;
assign img[13117] = 175;
assign img[13118] = 138;
assign img[13119] = 136;
assign img[13120] = 248;
assign img[13121] = 223;
assign img[13122] = 137;
assign img[13123] = 234;
assign img[13124] = 238;
assign img[13125] = 255;
assign img[13126] = 191;
assign img[13127] = 139;
assign img[13128] = 136;
assign img[13129] = 238;
assign img[13130] = 254;
assign img[13131] = 191;
assign img[13132] = 187;
assign img[13133] = 187;
assign img[13134] = 187;
assign img[13135] = 251;
assign img[13136] = 143;
assign img[13137] = 234;
assign img[13138] = 238;
assign img[13139] = 238;
assign img[13140] = 238;
assign img[13141] = 206;
assign img[13142] = 136;
assign img[13143] = 204;
assign img[13144] = 140;
assign img[13145] = 152;
assign img[13146] = 185;
assign img[13147] = 155;
assign img[13148] = 217;
assign img[13149] = 221;
assign img[13150] = 153;
assign img[13151] = 153;
assign img[13152] = 153;
assign img[13153] = 153;
assign img[13154] = 217;
assign img[13155] = 255;
assign img[13156] = 255;
assign img[13157] = 223;
assign img[13158] = 189;
assign img[13159] = 186;
assign img[13160] = 234;
assign img[13161] = 206;
assign img[13162] = 220;
assign img[13163] = 157;
assign img[13164] = 153;
assign img[13165] = 217;
assign img[13166] = 185;
assign img[13167] = 187;
assign img[13168] = 187;
assign img[13169] = 255;
assign img[13170] = 255;
assign img[13171] = 223;
assign img[13172] = 253;
assign img[13173] = 191;
assign img[13174] = 223;
assign img[13175] = 255;
assign img[13176] = 255;
assign img[13177] = 255;
assign img[13178] = 171;
assign img[13179] = 170;
assign img[13180] = 170;
assign img[13181] = 234;
assign img[13182] = 174;
assign img[13183] = 234;
assign img[13184] = 16;
assign img[13185] = 221;
assign img[13186] = 253;
assign img[13187] = 255;
assign img[13188] = 255;
assign img[13189] = 207;
assign img[13190] = 236;
assign img[13191] = 206;
assign img[13192] = 204;
assign img[13193] = 206;
assign img[13194] = 220;
assign img[13195] = 237;
assign img[13196] = 238;
assign img[13197] = 238;
assign img[13198] = 206;
assign img[13199] = 140;
assign img[13200] = 200;
assign img[13201] = 204;
assign img[13202] = 204;
assign img[13203] = 140;
assign img[13204] = 200;
assign img[13205] = 238;
assign img[13206] = 174;
assign img[13207] = 238;
assign img[13208] = 238;
assign img[13209] = 191;
assign img[13210] = 153;
assign img[13211] = 201;
assign img[13212] = 136;
assign img[13213] = 204;
assign img[13214] = 136;
assign img[13215] = 136;
assign img[13216] = 136;
assign img[13217] = 153;
assign img[13218] = 185;
assign img[13219] = 187;
assign img[13220] = 171;
assign img[13221] = 138;
assign img[13222] = 136;
assign img[13223] = 204;
assign img[13224] = 204;
assign img[13225] = 238;
assign img[13226] = 254;
assign img[13227] = 255;
assign img[13228] = 153;
assign img[13229] = 137;
assign img[13230] = 232;
assign img[13231] = 239;
assign img[13232] = 238;
assign img[13233] = 206;
assign img[13234] = 220;
assign img[13235] = 255;
assign img[13236] = 170;
assign img[13237] = 138;
assign img[13238] = 152;
assign img[13239] = 223;
assign img[13240] = 204;
assign img[13241] = 204;
assign img[13242] = 236;
assign img[13243] = 238;
assign img[13244] = 238;
assign img[13245] = 142;
assign img[13246] = 152;
assign img[13247] = 201;
assign img[13248] = 204;
assign img[13249] = 174;
assign img[13250] = 139;
assign img[13251] = 232;
assign img[13252] = 238;
assign img[13253] = 174;
assign img[13254] = 250;
assign img[13255] = 255;
assign img[13256] = 204;
assign img[13257] = 204;
assign img[13258] = 136;
assign img[13259] = 253;
assign img[13260] = 255;
assign img[13261] = 191;
assign img[13262] = 255;
assign img[13263] = 255;
assign img[13264] = 238;
assign img[13265] = 238;
assign img[13266] = 238;
assign img[13267] = 254;
assign img[13268] = 255;
assign img[13269] = 159;
assign img[13270] = 153;
assign img[13271] = 255;
assign img[13272] = 255;
assign img[13273] = 223;
assign img[13274] = 221;
assign img[13275] = 189;
assign img[13276] = 136;
assign img[13277] = 191;
assign img[13278] = 187;
assign img[13279] = 155;
assign img[13280] = 185;
assign img[13281] = 171;
assign img[13282] = 170;
assign img[13283] = 254;
assign img[13284] = 255;
assign img[13285] = 191;
assign img[13286] = 138;
assign img[13287] = 187;
assign img[13288] = 251;
assign img[13289] = 191;
assign img[13290] = 251;
assign img[13291] = 255;
assign img[13292] = 140;
assign img[13293] = 136;
assign img[13294] = 200;
assign img[13295] = 204;
assign img[13296] = 140;
assign img[13297] = 136;
assign img[13298] = 232;
assign img[13299] = 190;
assign img[13300] = 187;
assign img[13301] = 187;
assign img[13302] = 221;
assign img[13303] = 221;
assign img[13304] = 221;
assign img[13305] = 253;
assign img[13306] = 223;
assign img[13307] = 204;
assign img[13308] = 220;
assign img[13309] = 255;
assign img[13310] = 255;
assign img[13311] = 255;
assign img[13312] = 96;
assign img[13313] = 206;
assign img[13314] = 220;
assign img[13315] = 221;
assign img[13316] = 153;
assign img[13317] = 187;
assign img[13318] = 171;
assign img[13319] = 251;
assign img[13320] = 255;
assign img[13321] = 255;
assign img[13322] = 255;
assign img[13323] = 255;
assign img[13324] = 221;
assign img[13325] = 221;
assign img[13326] = 253;
assign img[13327] = 159;
assign img[13328] = 153;
assign img[13329] = 191;
assign img[13330] = 223;
assign img[13331] = 157;
assign img[13332] = 153;
assign img[13333] = 221;
assign img[13334] = 157;
assign img[13335] = 251;
assign img[13336] = 255;
assign img[13337] = 255;
assign img[13338] = 170;
assign img[13339] = 234;
assign img[13340] = 238;
assign img[13341] = 255;
assign img[13342] = 191;
assign img[13343] = 171;
assign img[13344] = 136;
assign img[13345] = 248;
assign img[13346] = 191;
assign img[13347] = 235;
assign img[13348] = 186;
assign img[13349] = 187;
assign img[13350] = 155;
assign img[13351] = 153;
assign img[13352] = 232;
assign img[13353] = 222;
assign img[13354] = 204;
assign img[13355] = 238;
assign img[13356] = 138;
assign img[13357] = 184;
assign img[13358] = 251;
assign img[13359] = 191;
assign img[13360] = 251;
assign img[13361] = 239;
assign img[13362] = 174;
assign img[13363] = 170;
assign img[13364] = 170;
assign img[13365] = 170;
assign img[13366] = 136;
assign img[13367] = 204;
assign img[13368] = 204;
assign img[13369] = 204;
assign img[13370] = 140;
assign img[13371] = 137;
assign img[13372] = 232;
assign img[13373] = 142;
assign img[13374] = 136;
assign img[13375] = 234;
assign img[13376] = 238;
assign img[13377] = 191;
assign img[13378] = 155;
assign img[13379] = 251;
assign img[13380] = 239;
assign img[13381] = 255;
assign img[13382] = 255;
assign img[13383] = 255;
assign img[13384] = 255;
assign img[13385] = 255;
assign img[13386] = 238;
assign img[13387] = 204;
assign img[13388] = 140;
assign img[13389] = 190;
assign img[13390] = 187;
assign img[13391] = 187;
assign img[13392] = 187;
assign img[13393] = 251;
assign img[13394] = 255;
assign img[13395] = 207;
assign img[13396] = 236;
assign img[13397] = 158;
assign img[13398] = 153;
assign img[13399] = 255;
assign img[13400] = 207;
assign img[13401] = 204;
assign img[13402] = 220;
assign img[13403] = 159;
assign img[13404] = 217;
assign img[13405] = 175;
assign img[13406] = 234;
assign img[13407] = 239;
assign img[13408] = 187;
assign img[13409] = 187;
assign img[13410] = 251;
assign img[13411] = 255;
assign img[13412] = 255;
assign img[13413] = 191;
assign img[13414] = 136;
assign img[13415] = 200;
assign img[13416] = 236;
assign img[13417] = 238;
assign img[13418] = 238;
assign img[13419] = 255;
assign img[13420] = 170;
assign img[13421] = 201;
assign img[13422] = 253;
assign img[13423] = 239;
assign img[13424] = 254;
assign img[13425] = 187;
assign img[13426] = 155;
assign img[13427] = 153;
assign img[13428] = 217;
assign img[13429] = 205;
assign img[13430] = 204;
assign img[13431] = 254;
assign img[13432] = 255;
assign img[13433] = 255;
assign img[13434] = 238;
assign img[13435] = 255;
assign img[13436] = 255;
assign img[13437] = 255;
assign img[13438] = 251;
assign img[13439] = 255;
assign img[13440] = 0;
assign img[13441] = 137;
assign img[13442] = 232;
assign img[13443] = 238;
assign img[13444] = 238;
assign img[13445] = 255;
assign img[13446] = 157;
assign img[13447] = 153;
assign img[13448] = 217;
assign img[13449] = 255;
assign img[13450] = 255;
assign img[13451] = 191;
assign img[13452] = 187;
assign img[13453] = 187;
assign img[13454] = 251;
assign img[13455] = 191;
assign img[13456] = 255;
assign img[13457] = 223;
assign img[13458] = 204;
assign img[13459] = 140;
assign img[13460] = 184;
assign img[13461] = 187;
assign img[13462] = 207;
assign img[13463] = 204;
assign img[13464] = 220;
assign img[13465] = 157;
assign img[13466] = 204;
assign img[13467] = 253;
assign img[13468] = 255;
assign img[13469] = 255;
assign img[13470] = 255;
assign img[13471] = 207;
assign img[13472] = 136;
assign img[13473] = 136;
assign img[13474] = 200;
assign img[13475] = 140;
assign img[13476] = 136;
assign img[13477] = 168;
assign img[13478] = 234;
assign img[13479] = 174;
assign img[13480] = 187;
assign img[13481] = 155;
assign img[13482] = 170;
assign img[13483] = 138;
assign img[13484] = 136;
assign img[13485] = 136;
assign img[13486] = 217;
assign img[13487] = 157;
assign img[13488] = 185;
assign img[13489] = 155;
assign img[13490] = 232;
assign img[13491] = 190;
assign img[13492] = 153;
assign img[13493] = 251;
assign img[13494] = 136;
assign img[13495] = 137;
assign img[13496] = 136;
assign img[13497] = 136;
assign img[13498] = 136;
assign img[13499] = 136;
assign img[13500] = 200;
assign img[13501] = 140;
assign img[13502] = 248;
assign img[13503] = 255;
assign img[13504] = 255;
assign img[13505] = 255;
assign img[13506] = 155;
assign img[13507] = 187;
assign img[13508] = 187;
assign img[13509] = 187;
assign img[13510] = 187;
assign img[13511] = 187;
assign img[13512] = 170;
assign img[13513] = 250;
assign img[13514] = 239;
assign img[13515] = 238;
assign img[13516] = 170;
assign img[13517] = 202;
assign img[13518] = 136;
assign img[13519] = 206;
assign img[13520] = 136;
assign img[13521] = 217;
assign img[13522] = 237;
assign img[13523] = 190;
assign img[13524] = 171;
assign img[13525] = 138;
assign img[13526] = 136;
assign img[13527] = 136;
assign img[13528] = 186;
assign img[13529] = 251;
assign img[13530] = 187;
assign img[13531] = 155;
assign img[13532] = 153;
assign img[13533] = 217;
assign img[13534] = 221;
assign img[13535] = 205;
assign img[13536] = 136;
assign img[13537] = 168;
assign img[13538] = 234;
assign img[13539] = 238;
assign img[13540] = 238;
assign img[13541] = 223;
assign img[13542] = 205;
assign img[13543] = 221;
assign img[13544] = 221;
assign img[13545] = 221;
assign img[13546] = 221;
assign img[13547] = 255;
assign img[13548] = 255;
assign img[13549] = 255;
assign img[13550] = 221;
assign img[13551] = 221;
assign img[13552] = 221;
assign img[13553] = 221;
assign img[13554] = 221;
assign img[13555] = 157;
assign img[13556] = 153;
assign img[13557] = 153;
assign img[13558] = 153;
assign img[13559] = 235;
assign img[13560] = 255;
assign img[13561] = 171;
assign img[13562] = 136;
assign img[13563] = 136;
assign img[13564] = 232;
assign img[13565] = 238;
assign img[13566] = 238;
assign img[13567] = 186;
assign img[13568] = 96;
assign img[13569] = 206;
assign img[13570] = 252;
assign img[13571] = 239;
assign img[13572] = 206;
assign img[13573] = 204;
assign img[13574] = 188;
assign img[13575] = 223;
assign img[13576] = 236;
assign img[13577] = 238;
assign img[13578] = 238;
assign img[13579] = 238;
assign img[13580] = 238;
assign img[13581] = 204;
assign img[13582] = 204;
assign img[13583] = 156;
assign img[13584] = 153;
assign img[13585] = 153;
assign img[13586] = 153;
assign img[13587] = 157;
assign img[13588] = 153;
assign img[13589] = 153;
assign img[13590] = 153;
assign img[13591] = 153;
assign img[13592] = 253;
assign img[13593] = 175;
assign img[13594] = 174;
assign img[13595] = 239;
assign img[13596] = 238;
assign img[13597] = 238;
assign img[13598] = 238;
assign img[13599] = 143;
assign img[13600] = 136;
assign img[13601] = 153;
assign img[13602] = 153;
assign img[13603] = 137;
assign img[13604] = 168;
assign img[13605] = 186;
assign img[13606] = 171;
assign img[13607] = 170;
assign img[13608] = 234;
assign img[13609] = 220;
assign img[13610] = 205;
assign img[13611] = 204;
assign img[13612] = 220;
assign img[13613] = 239;
assign img[13614] = 236;
assign img[13615] = 255;
assign img[13616] = 255;
assign img[13617] = 255;
assign img[13618] = 255;
assign img[13619] = 238;
assign img[13620] = 238;
assign img[13621] = 222;
assign img[13622] = 221;
assign img[13623] = 205;
assign img[13624] = 140;
assign img[13625] = 152;
assign img[13626] = 153;
assign img[13627] = 153;
assign img[13628] = 168;
assign img[13629] = 174;
assign img[13630] = 186;
assign img[13631] = 219;
assign img[13632] = 221;
assign img[13633] = 221;
assign img[13634] = 253;
assign img[13635] = 255;
assign img[13636] = 239;
assign img[13637] = 255;
assign img[13638] = 187;
assign img[13639] = 187;
assign img[13640] = 251;
assign img[13641] = 207;
assign img[13642] = 220;
assign img[13643] = 205;
assign img[13644] = 204;
assign img[13645] = 239;
assign img[13646] = 238;
assign img[13647] = 238;
assign img[13648] = 238;
assign img[13649] = 238;
assign img[13650] = 238;
assign img[13651] = 254;
assign img[13652] = 238;
assign img[13653] = 238;
assign img[13654] = 204;
assign img[13655] = 204;
assign img[13656] = 157;
assign img[13657] = 185;
assign img[13658] = 251;
assign img[13659] = 191;
assign img[13660] = 187;
assign img[13661] = 255;
assign img[13662] = 255;
assign img[13663] = 159;
assign img[13664] = 137;
assign img[13665] = 217;
assign img[13666] = 221;
assign img[13667] = 255;
assign img[13668] = 238;
assign img[13669] = 254;
assign img[13670] = 255;
assign img[13671] = 239;
assign img[13672] = 238;
assign img[13673] = 238;
assign img[13674] = 170;
assign img[13675] = 170;
assign img[13676] = 254;
assign img[13677] = 207;
assign img[13678] = 204;
assign img[13679] = 140;
assign img[13680] = 136;
assign img[13681] = 201;
assign img[13682] = 221;
assign img[13683] = 205;
assign img[13684] = 189;
assign img[13685] = 187;
assign img[13686] = 251;
assign img[13687] = 255;
assign img[13688] = 207;
assign img[13689] = 204;
assign img[13690] = 168;
assign img[13691] = 254;
assign img[13692] = 187;
assign img[13693] = 255;
assign img[13694] = 223;
assign img[13695] = 255;
assign img[13696] = 80;
assign img[13697] = 245;
assign img[13698] = 255;
assign img[13699] = 255;
assign img[13700] = 223;
assign img[13701] = 255;
assign img[13702] = 223;
assign img[13703] = 221;
assign img[13704] = 253;
assign img[13705] = 223;
assign img[13706] = 221;
assign img[13707] = 221;
assign img[13708] = 221;
assign img[13709] = 239;
assign img[13710] = 186;
assign img[13711] = 159;
assign img[13712] = 153;
assign img[13713] = 189;
assign img[13714] = 155;
assign img[13715] = 253;
assign img[13716] = 251;
assign img[13717] = 255;
assign img[13718] = 239;
assign img[13719] = 238;
assign img[13720] = 238;
assign img[13721] = 238;
assign img[13722] = 142;
assign img[13723] = 206;
assign img[13724] = 255;
assign img[13725] = 255;
assign img[13726] = 205;
assign img[13727] = 174;
assign img[13728] = 152;
assign img[13729] = 155;
assign img[13730] = 187;
assign img[13731] = 187;
assign img[13732] = 187;
assign img[13733] = 171;
assign img[13734] = 170;
assign img[13735] = 190;
assign img[13736] = 239;
assign img[13737] = 238;
assign img[13738] = 140;
assign img[13739] = 170;
assign img[13740] = 186;
assign img[13741] = 155;
assign img[13742] = 234;
assign img[13743] = 255;
assign img[13744] = 238;
assign img[13745] = 238;
assign img[13746] = 238;
assign img[13747] = 238;
assign img[13748] = 206;
assign img[13749] = 238;
assign img[13750] = 174;
assign img[13751] = 238;
assign img[13752] = 205;
assign img[13753] = 204;
assign img[13754] = 152;
assign img[13755] = 153;
assign img[13756] = 249;
assign img[13757] = 255;
assign img[13758] = 187;
assign img[13759] = 171;
assign img[13760] = 251;
assign img[13761] = 190;
assign img[13762] = 170;
assign img[13763] = 238;
assign img[13764] = 174;
assign img[13765] = 170;
assign img[13766] = 170;
assign img[13767] = 170;
assign img[13768] = 250;
assign img[13769] = 191;
assign img[13770] = 251;
assign img[13771] = 239;
assign img[13772] = 238;
assign img[13773] = 206;
assign img[13774] = 252;
assign img[13775] = 255;
assign img[13776] = 239;
assign img[13777] = 238;
assign img[13778] = 238;
assign img[13779] = 190;
assign img[13780] = 187;
assign img[13781] = 187;
assign img[13782] = 234;
assign img[13783] = 239;
assign img[13784] = 174;
assign img[13785] = 171;
assign img[13786] = 170;
assign img[13787] = 186;
assign img[13788] = 187;
assign img[13789] = 187;
assign img[13790] = 217;
assign img[13791] = 253;
assign img[13792] = 187;
assign img[13793] = 187;
assign img[13794] = 234;
assign img[13795] = 238;
assign img[13796] = 220;
assign img[13797] = 141;
assign img[13798] = 184;
assign img[13799] = 139;
assign img[13800] = 152;
assign img[13801] = 223;
assign img[13802] = 236;
assign img[13803] = 238;
assign img[13804] = 238;
assign img[13805] = 238;
assign img[13806] = 254;
assign img[13807] = 255;
assign img[13808] = 191;
assign img[13809] = 221;
assign img[13810] = 237;
assign img[13811] = 255;
assign img[13812] = 255;
assign img[13813] = 239;
assign img[13814] = 254;
assign img[13815] = 255;
assign img[13816] = 255;
assign img[13817] = 223;
assign img[13818] = 255;
assign img[13819] = 223;
assign img[13820] = 221;
assign img[13821] = 253;
assign img[13822] = 255;
assign img[13823] = 255;
assign img[13824] = 96;
assign img[13825] = 238;
assign img[13826] = 254;
assign img[13827] = 255;
assign img[13828] = 238;
assign img[13829] = 238;
assign img[13830] = 174;
assign img[13831] = 254;
assign img[13832] = 255;
assign img[13833] = 255;
assign img[13834] = 238;
assign img[13835] = 238;
assign img[13836] = 170;
assign img[13837] = 238;
assign img[13838] = 238;
assign img[13839] = 174;
assign img[13840] = 170;
assign img[13841] = 154;
assign img[13842] = 153;
assign img[13843] = 185;
assign img[13844] = 155;
assign img[13845] = 157;
assign img[13846] = 205;
assign img[13847] = 204;
assign img[13848] = 204;
assign img[13849] = 204;
assign img[13850] = 236;
assign img[13851] = 238;
assign img[13852] = 238;
assign img[13853] = 238;
assign img[13854] = 206;
assign img[13855] = 140;
assign img[13856] = 136;
assign img[13857] = 200;
assign img[13858] = 204;
assign img[13859] = 254;
assign img[13860] = 191;
assign img[13861] = 155;
assign img[13862] = 137;
assign img[13863] = 140;
assign img[13864] = 220;
assign img[13865] = 237;
assign img[13866] = 238;
assign img[13867] = 238;
assign img[13868] = 238;
assign img[13869] = 207;
assign img[13870] = 236;
assign img[13871] = 174;
assign img[13872] = 238;
assign img[13873] = 239;
assign img[13874] = 238;
assign img[13875] = 175;
assign img[13876] = 187;
assign img[13877] = 251;
assign img[13878] = 239;
assign img[13879] = 223;
assign img[13880] = 253;
assign img[13881] = 255;
assign img[13882] = 221;
assign img[13883] = 253;
assign img[13884] = 239;
assign img[13885] = 206;
assign img[13886] = 236;
assign img[13887] = 238;
assign img[13888] = 204;
assign img[13889] = 252;
assign img[13890] = 223;
assign img[13891] = 237;
assign img[13892] = 254;
assign img[13893] = 255;
assign img[13894] = 221;
assign img[13895] = 223;
assign img[13896] = 255;
assign img[13897] = 221;
assign img[13898] = 253;
assign img[13899] = 191;
assign img[13900] = 187;
assign img[13901] = 187;
assign img[13902] = 187;
assign img[13903] = 255;
assign img[13904] = 255;
assign img[13905] = 255;
assign img[13906] = 239;
assign img[13907] = 238;
assign img[13908] = 254;
assign img[13909] = 239;
assign img[13910] = 170;
assign img[13911] = 206;
assign img[13912] = 236;
assign img[13913] = 238;
assign img[13914] = 222;
assign img[13915] = 157;
assign img[13916] = 249;
assign img[13917] = 223;
assign img[13918] = 253;
assign img[13919] = 191;
assign img[13920] = 138;
assign img[13921] = 200;
assign img[13922] = 204;
assign img[13923] = 206;
assign img[13924] = 204;
assign img[13925] = 236;
assign img[13926] = 238;
assign img[13927] = 238;
assign img[13928] = 254;
assign img[13929] = 223;
assign img[13930] = 204;
assign img[13931] = 204;
assign img[13932] = 204;
assign img[13933] = 206;
assign img[13934] = 204;
assign img[13935] = 236;
assign img[13936] = 170;
assign img[13937] = 186;
assign img[13938] = 219;
assign img[13939] = 221;
assign img[13940] = 221;
assign img[13941] = 191;
assign img[13942] = 171;
assign img[13943] = 238;
assign img[13944] = 238;
assign img[13945] = 191;
assign img[13946] = 255;
assign img[13947] = 175;
assign img[13948] = 170;
assign img[13949] = 254;
assign img[13950] = 255;
assign img[13951] = 255;
assign img[13952] = 96;
assign img[13953] = 238;
assign img[13954] = 254;
assign img[13955] = 255;
assign img[13956] = 255;
assign img[13957] = 255;
assign img[13958] = 153;
assign img[13959] = 251;
assign img[13960] = 255;
assign img[13961] = 255;
assign img[13962] = 238;
assign img[13963] = 204;
assign img[13964] = 140;
assign img[13965] = 169;
assign img[13966] = 155;
assign img[13967] = 153;
assign img[13968] = 137;
assign img[13969] = 170;
assign img[13970] = 234;
assign img[13971] = 174;
assign img[13972] = 202;
assign img[13973] = 238;
assign img[13974] = 206;
assign img[13975] = 204;
assign img[13976] = 204;
assign img[13977] = 206;
assign img[13978] = 136;
assign img[13979] = 234;
assign img[13980] = 238;
assign img[13981] = 238;
assign img[13982] = 190;
assign img[13983] = 191;
assign img[13984] = 187;
assign img[13985] = 251;
assign img[13986] = 207;
assign img[13987] = 220;
assign img[13988] = 221;
assign img[13989] = 221;
assign img[13990] = 221;
assign img[13991] = 205;
assign img[13992] = 221;
assign img[13993] = 221;
assign img[13994] = 223;
assign img[13995] = 140;
assign img[13996] = 236;
assign img[13997] = 174;
assign img[13998] = 186;
assign img[13999] = 191;
assign img[14000] = 170;
assign img[14001] = 138;
assign img[14002] = 200;
assign img[14003] = 204;
assign img[14004] = 156;
assign img[14005] = 153;
assign img[14006] = 153;
assign img[14007] = 137;
assign img[14008] = 168;
assign img[14009] = 239;
assign img[14010] = 255;
assign img[14011] = 255;
assign img[14012] = 255;
assign img[14013] = 191;
assign img[14014] = 155;
assign img[14015] = 255;
assign img[14016] = 255;
assign img[14017] = 239;
assign img[14018] = 238;
assign img[14019] = 238;
assign img[14020] = 238;
assign img[14021] = 238;
assign img[14022] = 136;
assign img[14023] = 220;
assign img[14024] = 153;
assign img[14025] = 153;
assign img[14026] = 153;
assign img[14027] = 153;
assign img[14028] = 153;
assign img[14029] = 204;
assign img[14030] = 204;
assign img[14031] = 238;
assign img[14032] = 174;
assign img[14033] = 170;
assign img[14034] = 186;
assign img[14035] = 187;
assign img[14036] = 187;
assign img[14037] = 171;
assign img[14038] = 234;
assign img[14039] = 238;
assign img[14040] = 204;
assign img[14041] = 238;
assign img[14042] = 238;
assign img[14043] = 142;
assign img[14044] = 204;
assign img[14045] = 204;
assign img[14046] = 236;
assign img[14047] = 238;
assign img[14048] = 238;
assign img[14049] = 238;
assign img[14050] = 238;
assign img[14051] = 238;
assign img[14052] = 238;
assign img[14053] = 174;
assign img[14054] = 254;
assign img[14055] = 255;
assign img[14056] = 255;
assign img[14057] = 223;
assign img[14058] = 253;
assign img[14059] = 239;
assign img[14060] = 204;
assign img[14061] = 238;
assign img[14062] = 238;
assign img[14063] = 238;
assign img[14064] = 254;
assign img[14065] = 191;
assign img[14066] = 171;
assign img[14067] = 154;
assign img[14068] = 217;
assign img[14069] = 205;
assign img[14070] = 204;
assign img[14071] = 236;
assign img[14072] = 238;
assign img[14073] = 174;
assign img[14074] = 186;
assign img[14075] = 191;
assign img[14076] = 187;
assign img[14077] = 251;
assign img[14078] = 255;
assign img[14079] = 255;
assign img[14080] = 96;
assign img[14081] = 223;
assign img[14082] = 253;
assign img[14083] = 239;
assign img[14084] = 154;
assign img[14085] = 205;
assign img[14086] = 204;
assign img[14087] = 252;
assign img[14088] = 254;
assign img[14089] = 255;
assign img[14090] = 191;
assign img[14091] = 155;
assign img[14092] = 153;
assign img[14093] = 200;
assign img[14094] = 220;
assign img[14095] = 141;
assign img[14096] = 204;
assign img[14097] = 204;
assign img[14098] = 204;
assign img[14099] = 254;
assign img[14100] = 255;
assign img[14101] = 191;
assign img[14102] = 187;
assign img[14103] = 251;
assign img[14104] = 255;
assign img[14105] = 223;
assign img[14106] = 221;
assign img[14107] = 221;
assign img[14108] = 253;
assign img[14109] = 223;
assign img[14110] = 253;
assign img[14111] = 138;
assign img[14112] = 136;
assign img[14113] = 232;
assign img[14114] = 238;
assign img[14115] = 238;
assign img[14116] = 255;
assign img[14117] = 191;
assign img[14118] = 187;
assign img[14119] = 187;
assign img[14120] = 136;
assign img[14121] = 170;
assign img[14122] = 136;
assign img[14123] = 136;
assign img[14124] = 136;
assign img[14125] = 156;
assign img[14126] = 253;
assign img[14127] = 191;
assign img[14128] = 187;
assign img[14129] = 187;
assign img[14130] = 170;
assign img[14131] = 170;
assign img[14132] = 155;
assign img[14133] = 251;
assign img[14134] = 239;
assign img[14135] = 238;
assign img[14136] = 206;
assign img[14137] = 204;
assign img[14138] = 136;
assign img[14139] = 232;
assign img[14140] = 190;
assign img[14141] = 155;
assign img[14142] = 153;
assign img[14143] = 253;
assign img[14144] = 238;
assign img[14145] = 254;
assign img[14146] = 153;
assign img[14147] = 153;
assign img[14148] = 249;
assign img[14149] = 191;
assign img[14150] = 153;
assign img[14151] = 255;
assign img[14152] = 255;
assign img[14153] = 223;
assign img[14154] = 238;
assign img[14155] = 142;
assign img[14156] = 136;
assign img[14157] = 153;
assign img[14158] = 137;
assign img[14159] = 170;
assign img[14160] = 154;
assign img[14161] = 251;
assign img[14162] = 239;
assign img[14163] = 206;
assign img[14164] = 204;
assign img[14165] = 172;
assign img[14166] = 138;
assign img[14167] = 253;
assign img[14168] = 159;
assign img[14169] = 137;
assign img[14170] = 136;
assign img[14171] = 136;
assign img[14172] = 232;
assign img[14173] = 238;
assign img[14174] = 238;
assign img[14175] = 206;
assign img[14176] = 204;
assign img[14177] = 238;
assign img[14178] = 170;
assign img[14179] = 238;
assign img[14180] = 206;
assign img[14181] = 238;
assign img[14182] = 222;
assign img[14183] = 221;
assign img[14184] = 255;
assign img[14185] = 255;
assign img[14186] = 255;
assign img[14187] = 255;
assign img[14188] = 171;
assign img[14189] = 234;
assign img[14190] = 238;
assign img[14191] = 238;
assign img[14192] = 140;
assign img[14193] = 238;
assign img[14194] = 238;
assign img[14195] = 140;
assign img[14196] = 170;
assign img[14197] = 170;
assign img[14198] = 234;
assign img[14199] = 238;
assign img[14200] = 238;
assign img[14201] = 238;
assign img[14202] = 204;
assign img[14203] = 204;
assign img[14204] = 236;
assign img[14205] = 255;
assign img[14206] = 207;
assign img[14207] = 236;
assign img[14208] = 96;
assign img[14209] = 206;
assign img[14210] = 204;
assign img[14211] = 221;
assign img[14212] = 221;
assign img[14213] = 221;
assign img[14214] = 221;
assign img[14215] = 223;
assign img[14216] = 221;
assign img[14217] = 207;
assign img[14218] = 204;
assign img[14219] = 140;
assign img[14220] = 152;
assign img[14221] = 169;
assign img[14222] = 250;
assign img[14223] = 255;
assign img[14224] = 255;
assign img[14225] = 191;
assign img[14226] = 255;
assign img[14227] = 255;
assign img[14228] = 171;
assign img[14229] = 239;
assign img[14230] = 238;
assign img[14231] = 238;
assign img[14232] = 238;
assign img[14233] = 238;
assign img[14234] = 238;
assign img[14235] = 254;
assign img[14236] = 221;
assign img[14237] = 255;
assign img[14238] = 238;
assign img[14239] = 142;
assign img[14240] = 136;
assign img[14241] = 200;
assign img[14242] = 204;
assign img[14243] = 220;
assign img[14244] = 221;
assign img[14245] = 255;
assign img[14246] = 204;
assign img[14247] = 238;
assign img[14248] = 254;
assign img[14249] = 255;
assign img[14250] = 187;
assign img[14251] = 187;
assign img[14252] = 187;
assign img[14253] = 187;
assign img[14254] = 251;
assign img[14255] = 255;
assign img[14256] = 238;
assign img[14257] = 238;
assign img[14258] = 255;
assign img[14259] = 174;
assign img[14260] = 138;
assign img[14261] = 136;
assign img[14262] = 184;
assign img[14263] = 171;
assign img[14264] = 218;
assign img[14265] = 221;
assign img[14266] = 221;
assign img[14267] = 153;
assign img[14268] = 232;
assign img[14269] = 223;
assign img[14270] = 153;
assign img[14271] = 221;
assign img[14272] = 221;
assign img[14273] = 239;
assign img[14274] = 204;
assign img[14275] = 221;
assign img[14276] = 141;
assign img[14277] = 140;
assign img[14278] = 170;
assign img[14279] = 204;
assign img[14280] = 204;
assign img[14281] = 174;
assign img[14282] = 138;
assign img[14283] = 136;
assign img[14284] = 184;
assign img[14285] = 235;
assign img[14286] = 238;
assign img[14287] = 238;
assign img[14288] = 206;
assign img[14289] = 238;
assign img[14290] = 206;
assign img[14291] = 140;
assign img[14292] = 184;
assign img[14293] = 187;
assign img[14294] = 187;
assign img[14295] = 251;
assign img[14296] = 255;
assign img[14297] = 239;
assign img[14298] = 206;
assign img[14299] = 204;
assign img[14300] = 236;
assign img[14301] = 207;
assign img[14302] = 221;
assign img[14303] = 157;
assign img[14304] = 153;
assign img[14305] = 153;
assign img[14306] = 201;
assign img[14307] = 255;
assign img[14308] = 255;
assign img[14309] = 255;
assign img[14310] = 223;
assign img[14311] = 255;
assign img[14312] = 255;
assign img[14313] = 255;
assign img[14314] = 255;
assign img[14315] = 223;
assign img[14316] = 204;
assign img[14317] = 238;
assign img[14318] = 174;
assign img[14319] = 187;
assign img[14320] = 235;
assign img[14321] = 238;
assign img[14322] = 238;
assign img[14323] = 206;
assign img[14324] = 140;
assign img[14325] = 136;
assign img[14326] = 136;
assign img[14327] = 204;
assign img[14328] = 204;
assign img[14329] = 236;
assign img[14330] = 138;
assign img[14331] = 253;
assign img[14332] = 223;
assign img[14333] = 221;
assign img[14334] = 221;
assign img[14335] = 253;
assign img[14336] = 96;
assign img[14337] = 238;
assign img[14338] = 254;
assign img[14339] = 207;
assign img[14340] = 238;
assign img[14341] = 170;
assign img[14342] = 170;
assign img[14343] = 234;
assign img[14344] = 238;
assign img[14345] = 255;
assign img[14346] = 255;
assign img[14347] = 255;
assign img[14348] = 255;
assign img[14349] = 255;
assign img[14350] = 239;
assign img[14351] = 174;
assign img[14352] = 170;
assign img[14353] = 187;
assign img[14354] = 251;
assign img[14355] = 255;
assign img[14356] = 187;
assign img[14357] = 255;
assign img[14358] = 191;
assign img[14359] = 255;
assign img[14360] = 221;
assign img[14361] = 159;
assign img[14362] = 185;
assign img[14363] = 251;
assign img[14364] = 255;
assign img[14365] = 255;
assign img[14366] = 137;
assign img[14367] = 187;
assign img[14368] = 137;
assign img[14369] = 234;
assign img[14370] = 254;
assign img[14371] = 239;
assign img[14372] = 138;
assign img[14373] = 217;
assign img[14374] = 253;
assign img[14375] = 255;
assign img[14376] = 221;
assign img[14377] = 255;
assign img[14378] = 159;
assign img[14379] = 138;
assign img[14380] = 234;
assign img[14381] = 220;
assign img[14382] = 221;
assign img[14383] = 221;
assign img[14384] = 221;
assign img[14385] = 255;
assign img[14386] = 238;
assign img[14387] = 191;
assign img[14388] = 187;
assign img[14389] = 251;
assign img[14390] = 251;
assign img[14391] = 255;
assign img[14392] = 138;
assign img[14393] = 136;
assign img[14394] = 136;
assign img[14395] = 136;
assign img[14396] = 136;
assign img[14397] = 174;
assign img[14398] = 254;
assign img[14399] = 255;
assign img[14400] = 255;
assign img[14401] = 223;
assign img[14402] = 253;
assign img[14403] = 238;
assign img[14404] = 136;
assign img[14405] = 136;
assign img[14406] = 136;
assign img[14407] = 204;
assign img[14408] = 236;
assign img[14409] = 238;
assign img[14410] = 238;
assign img[14411] = 174;
assign img[14412] = 170;
assign img[14413] = 251;
assign img[14414] = 153;
assign img[14415] = 221;
assign img[14416] = 221;
assign img[14417] = 221;
assign img[14418] = 221;
assign img[14419] = 221;
assign img[14420] = 140;
assign img[14421] = 136;
assign img[14422] = 136;
assign img[14423] = 204;
assign img[14424] = 204;
assign img[14425] = 140;
assign img[14426] = 216;
assign img[14427] = 221;
assign img[14428] = 153;
assign img[14429] = 153;
assign img[14430] = 255;
assign img[14431] = 191;
assign img[14432] = 170;
assign img[14433] = 187;
assign img[14434] = 170;
assign img[14435] = 187;
assign img[14436] = 255;
assign img[14437] = 191;
assign img[14438] = 187;
assign img[14439] = 251;
assign img[14440] = 255;
assign img[14441] = 255;
assign img[14442] = 255;
assign img[14443] = 255;
assign img[14444] = 255;
assign img[14445] = 255;
assign img[14446] = 223;
assign img[14447] = 157;
assign img[14448] = 153;
assign img[14449] = 251;
assign img[14450] = 238;
assign img[14451] = 206;
assign img[14452] = 172;
assign img[14453] = 174;
assign img[14454] = 138;
assign img[14455] = 238;
assign img[14456] = 238;
assign img[14457] = 255;
assign img[14458] = 187;
assign img[14459] = 187;
assign img[14460] = 155;
assign img[14461] = 255;
assign img[14462] = 255;
assign img[14463] = 255;
assign img[14464] = 96;
assign img[14465] = 206;
assign img[14466] = 236;
assign img[14467] = 255;
assign img[14468] = 255;
assign img[14469] = 238;
assign img[14470] = 255;
assign img[14471] = 255;
assign img[14472] = 255;
assign img[14473] = 255;
assign img[14474] = 239;
assign img[14475] = 238;
assign img[14476] = 138;
assign img[14477] = 234;
assign img[14478] = 238;
assign img[14479] = 238;
assign img[14480] = 238;
assign img[14481] = 238;
assign img[14482] = 238;
assign img[14483] = 255;
assign img[14484] = 205;
assign img[14485] = 204;
assign img[14486] = 204;
assign img[14487] = 204;
assign img[14488] = 236;
assign img[14489] = 238;
assign img[14490] = 204;
assign img[14491] = 204;
assign img[14492] = 204;
assign img[14493] = 221;
assign img[14494] = 221;
assign img[14495] = 141;
assign img[14496] = 136;
assign img[14497] = 236;
assign img[14498] = 174;
assign img[14499] = 171;
assign img[14500] = 187;
assign img[14501] = 187;
assign img[14502] = 187;
assign img[14503] = 187;
assign img[14504] = 251;
assign img[14505] = 255;
assign img[14506] = 157;
assign img[14507] = 187;
assign img[14508] = 187;
assign img[14509] = 187;
assign img[14510] = 251;
assign img[14511] = 255;
assign img[14512] = 255;
assign img[14513] = 255;
assign img[14514] = 238;
assign img[14515] = 238;
assign img[14516] = 186;
assign img[14517] = 171;
assign img[14518] = 186;
assign img[14519] = 187;
assign img[14520] = 187;
assign img[14521] = 187;
assign img[14522] = 171;
assign img[14523] = 136;
assign img[14524] = 136;
assign img[14525] = 137;
assign img[14526] = 137;
assign img[14527] = 136;
assign img[14528] = 152;
assign img[14529] = 171;
assign img[14530] = 170;
assign img[14531] = 234;
assign img[14532] = 206;
assign img[14533] = 204;
assign img[14534] = 136;
assign img[14535] = 170;
assign img[14536] = 202;
assign img[14537] = 204;
assign img[14538] = 204;
assign img[14539] = 254;
assign img[14540] = 255;
assign img[14541] = 239;
assign img[14542] = 204;
assign img[14543] = 238;
assign img[14544] = 254;
assign img[14545] = 255;
assign img[14546] = 255;
assign img[14547] = 255;
assign img[14548] = 171;
assign img[14549] = 170;
assign img[14550] = 250;
assign img[14551] = 255;
assign img[14552] = 255;
assign img[14553] = 207;
assign img[14554] = 156;
assign img[14555] = 153;
assign img[14556] = 201;
assign img[14557] = 156;
assign img[14558] = 249;
assign img[14559] = 255;
assign img[14560] = 153;
assign img[14561] = 153;
assign img[14562] = 217;
assign img[14563] = 221;
assign img[14564] = 221;
assign img[14565] = 221;
assign img[14566] = 221;
assign img[14567] = 253;
assign img[14568] = 255;
assign img[14569] = 255;
assign img[14570] = 204;
assign img[14571] = 204;
assign img[14572] = 204;
assign img[14573] = 236;
assign img[14574] = 238;
assign img[14575] = 238;
assign img[14576] = 206;
assign img[14577] = 238;
assign img[14578] = 254;
assign img[14579] = 255;
assign img[14580] = 255;
assign img[14581] = 255;
assign img[14582] = 238;
assign img[14583] = 238;
assign img[14584] = 238;
assign img[14585] = 238;
assign img[14586] = 255;
assign img[14587] = 239;
assign img[14588] = 206;
assign img[14589] = 238;
assign img[14590] = 254;
assign img[14591] = 255;
assign img[14592] = 16;
assign img[14593] = 153;
assign img[14594] = 249;
assign img[14595] = 191;
assign img[14596] = 235;
assign img[14597] = 238;
assign img[14598] = 174;
assign img[14599] = 238;
assign img[14600] = 238;
assign img[14601] = 255;
assign img[14602] = 239;
assign img[14603] = 238;
assign img[14604] = 238;
assign img[14605] = 223;
assign img[14606] = 205;
assign img[14607] = 188;
assign img[14608] = 137;
assign img[14609] = 236;
assign img[14610] = 238;
assign img[14611] = 255;
assign img[14612] = 254;
assign img[14613] = 255;
assign img[14614] = 159;
assign img[14615] = 221;
assign img[14616] = 221;
assign img[14617] = 221;
assign img[14618] = 238;
assign img[14619] = 254;
assign img[14620] = 255;
assign img[14621] = 255;
assign img[14622] = 255;
assign img[14623] = 207;
assign img[14624] = 136;
assign img[14625] = 200;
assign img[14626] = 168;
assign img[14627] = 251;
assign img[14628] = 255;
assign img[14629] = 191;
assign img[14630] = 171;
assign img[14631] = 170;
assign img[14632] = 234;
assign img[14633] = 239;
assign img[14634] = 238;
assign img[14635] = 238;
assign img[14636] = 254;
assign img[14637] = 191;
assign img[14638] = 251;
assign img[14639] = 191;
assign img[14640] = 251;
assign img[14641] = 255;
assign img[14642] = 255;
assign img[14643] = 221;
assign img[14644] = 221;
assign img[14645] = 255;
assign img[14646] = 255;
assign img[14647] = 223;
assign img[14648] = 221;
assign img[14649] = 255;
assign img[14650] = 238;
assign img[14651] = 238;
assign img[14652] = 155;
assign img[14653] = 137;
assign img[14654] = 152;
assign img[14655] = 251;
assign img[14656] = 255;
assign img[14657] = 255;
assign img[14658] = 187;
assign img[14659] = 155;
assign img[14660] = 185;
assign img[14661] = 187;
assign img[14662] = 171;
assign img[14663] = 170;
assign img[14664] = 186;
assign img[14665] = 187;
assign img[14666] = 187;
assign img[14667] = 239;
assign img[14668] = 170;
assign img[14669] = 238;
assign img[14670] = 254;
assign img[14671] = 255;
assign img[14672] = 255;
assign img[14673] = 255;
assign img[14674] = 238;
assign img[14675] = 255;
assign img[14676] = 223;
assign img[14677] = 205;
assign img[14678] = 136;
assign img[14679] = 236;
assign img[14680] = 174;
assign img[14681] = 170;
assign img[14682] = 170;
assign img[14683] = 170;
assign img[14684] = 138;
assign img[14685] = 152;
assign img[14686] = 217;
assign img[14687] = 157;
assign img[14688] = 153;
assign img[14689] = 185;
assign img[14690] = 255;
assign img[14691] = 255;
assign img[14692] = 255;
assign img[14693] = 255;
assign img[14694] = 139;
assign img[14695] = 238;
assign img[14696] = 206;
assign img[14697] = 204;
assign img[14698] = 236;
assign img[14699] = 238;
assign img[14700] = 238;
assign img[14701] = 238;
assign img[14702] = 238;
assign img[14703] = 207;
assign img[14704] = 204;
assign img[14705] = 205;
assign img[14706] = 221;
assign img[14707] = 221;
assign img[14708] = 205;
assign img[14709] = 204;
assign img[14710] = 204;
assign img[14711] = 236;
assign img[14712] = 238;
assign img[14713] = 238;
assign img[14714] = 238;
assign img[14715] = 238;
assign img[14716] = 254;
assign img[14717] = 255;
assign img[14718] = 255;
assign img[14719] = 255;
assign img[14720] = 80;
assign img[14721] = 253;
assign img[14722] = 255;
assign img[14723] = 255;
assign img[14724] = 221;
assign img[14725] = 221;
assign img[14726] = 157;
assign img[14727] = 255;
assign img[14728] = 255;
assign img[14729] = 255;
assign img[14730] = 255;
assign img[14731] = 255;
assign img[14732] = 187;
assign img[14733] = 187;
assign img[14734] = 217;
assign img[14735] = 253;
assign img[14736] = 255;
assign img[14737] = 255;
assign img[14738] = 170;
assign img[14739] = 187;
assign img[14740] = 251;
assign img[14741] = 255;
assign img[14742] = 255;
assign img[14743] = 255;
assign img[14744] = 255;
assign img[14745] = 207;
assign img[14746] = 220;
assign img[14747] = 221;
assign img[14748] = 204;
assign img[14749] = 236;
assign img[14750] = 238;
assign img[14751] = 142;
assign img[14752] = 152;
assign img[14753] = 251;
assign img[14754] = 191;
assign img[14755] = 251;
assign img[14756] = 255;
assign img[14757] = 187;
assign img[14758] = 155;
assign img[14759] = 153;
assign img[14760] = 153;
assign img[14761] = 187;
assign img[14762] = 153;
assign img[14763] = 169;
assign img[14764] = 170;
assign img[14765] = 234;
assign img[14766] = 238;
assign img[14767] = 174;
assign img[14768] = 186;
assign img[14769] = 187;
assign img[14770] = 251;
assign img[14771] = 191;
assign img[14772] = 171;
assign img[14773] = 255;
assign img[14774] = 205;
assign img[14775] = 204;
assign img[14776] = 204;
assign img[14777] = 204;
assign img[14778] = 204;
assign img[14779] = 136;
assign img[14780] = 236;
assign img[14781] = 174;
assign img[14782] = 186;
assign img[14783] = 187;
assign img[14784] = 170;
assign img[14785] = 170;
assign img[14786] = 170;
assign img[14787] = 234;
assign img[14788] = 238;
assign img[14789] = 222;
assign img[14790] = 221;
assign img[14791] = 157;
assign img[14792] = 153;
assign img[14793] = 205;
assign img[14794] = 236;
assign img[14795] = 205;
assign img[14796] = 253;
assign img[14797] = 223;
assign img[14798] = 221;
assign img[14799] = 253;
assign img[14800] = 191;
assign img[14801] = 255;
assign img[14802] = 239;
assign img[14803] = 174;
assign img[14804] = 170;
assign img[14805] = 186;
assign img[14806] = 153;
assign img[14807] = 253;
assign img[14808] = 191;
assign img[14809] = 187;
assign img[14810] = 153;
assign img[14811] = 137;
assign img[14812] = 184;
assign img[14813] = 187;
assign img[14814] = 251;
assign img[14815] = 223;
assign img[14816] = 221;
assign img[14817] = 239;
assign img[14818] = 238;
assign img[14819] = 239;
assign img[14820] = 238;
assign img[14821] = 222;
assign img[14822] = 221;
assign img[14823] = 253;
assign img[14824] = 254;
assign img[14825] = 255;
assign img[14826] = 255;
assign img[14827] = 255;
assign img[14828] = 221;
assign img[14829] = 255;
assign img[14830] = 255;
assign img[14831] = 255;
assign img[14832] = 205;
assign img[14833] = 204;
assign img[14834] = 236;
assign img[14835] = 191;
assign img[14836] = 255;
assign img[14837] = 255;
assign img[14838] = 255;
assign img[14839] = 255;
assign img[14840] = 254;
assign img[14841] = 255;
assign img[14842] = 255;
assign img[14843] = 223;
assign img[14844] = 221;
assign img[14845] = 255;
assign img[14846] = 223;
assign img[14847] = 221;
assign img[14848] = 32;
assign img[14849] = 238;
assign img[14850] = 238;
assign img[14851] = 255;
assign img[14852] = 255;
assign img[14853] = 239;
assign img[14854] = 238;
assign img[14855] = 238;
assign img[14856] = 238;
assign img[14857] = 207;
assign img[14858] = 238;
assign img[14859] = 174;
assign img[14860] = 234;
assign img[14861] = 254;
assign img[14862] = 191;
assign img[14863] = 187;
assign img[14864] = 170;
assign img[14865] = 238;
assign img[14866] = 238;
assign img[14867] = 175;
assign img[14868] = 255;
assign img[14869] = 190;
assign img[14870] = 239;
assign img[14871] = 238;
assign img[14872] = 142;
assign img[14873] = 153;
assign img[14874] = 153;
assign img[14875] = 253;
assign img[14876] = 207;
assign img[14877] = 204;
assign img[14878] = 220;
assign img[14879] = 153;
assign img[14880] = 136;
assign img[14881] = 232;
assign img[14882] = 174;
assign img[14883] = 170;
assign img[14884] = 136;
assign img[14885] = 187;
assign img[14886] = 155;
assign img[14887] = 255;
assign img[14888] = 255;
assign img[14889] = 255;
assign img[14890] = 157;
assign img[14891] = 221;
assign img[14892] = 255;
assign img[14893] = 221;
assign img[14894] = 255;
assign img[14895] = 255;
assign img[14896] = 187;
assign img[14897] = 255;
assign img[14898] = 223;
assign img[14899] = 255;
assign img[14900] = 187;
assign img[14901] = 251;
assign img[14902] = 153;
assign img[14903] = 187;
assign img[14904] = 234;
assign img[14905] = 206;
assign img[14906] = 220;
assign img[14907] = 255;
assign img[14908] = 238;
assign img[14909] = 159;
assign img[14910] = 153;
assign img[14911] = 153;
assign img[14912] = 249;
assign img[14913] = 223;
assign img[14914] = 157;
assign img[14915] = 185;
assign img[14916] = 171;
assign img[14917] = 170;
assign img[14918] = 138;
assign img[14919] = 220;
assign img[14920] = 189;
assign img[14921] = 187;
assign img[14922] = 219;
assign img[14923] = 191;
assign img[14924] = 187;
assign img[14925] = 238;
assign img[14926] = 238;
assign img[14927] = 238;
assign img[14928] = 170;
assign img[14929] = 234;
assign img[14930] = 238;
assign img[14931] = 238;
assign img[14932] = 220;
assign img[14933] = 237;
assign img[14934] = 238;
assign img[14935] = 238;
assign img[14936] = 174;
assign img[14937] = 170;
assign img[14938] = 136;
assign img[14939] = 153;
assign img[14940] = 153;
assign img[14941] = 153;
assign img[14942] = 249;
assign img[14943] = 255;
assign img[14944] = 137;
assign img[14945] = 136;
assign img[14946] = 216;
assign img[14947] = 221;
assign img[14948] = 236;
assign img[14949] = 238;
assign img[14950] = 174;
assign img[14951] = 187;
assign img[14952] = 251;
assign img[14953] = 239;
assign img[14954] = 174;
assign img[14955] = 238;
assign img[14956] = 238;
assign img[14957] = 238;
assign img[14958] = 238;
assign img[14959] = 238;
assign img[14960] = 238;
assign img[14961] = 174;
assign img[14962] = 170;
assign img[14963] = 239;
assign img[14964] = 174;
assign img[14965] = 170;
assign img[14966] = 138;
assign img[14967] = 238;
assign img[14968] = 238;
assign img[14969] = 255;
assign img[14970] = 238;
assign img[14971] = 238;
assign img[14972] = 204;
assign img[14973] = 236;
assign img[14974] = 254;
assign img[14975] = 255;
assign img[14976] = 96;
assign img[14977] = 142;
assign img[14978] = 232;
assign img[14979] = 223;
assign img[14980] = 157;
assign img[14981] = 221;
assign img[14982] = 221;
assign img[14983] = 255;
assign img[14984] = 255;
assign img[14985] = 255;
assign img[14986] = 239;
assign img[14987] = 255;
assign img[14988] = 255;
assign img[14989] = 239;
assign img[14990] = 238;
assign img[14991] = 238;
assign img[14992] = 254;
assign img[14993] = 239;
assign img[14994] = 238;
assign img[14995] = 238;
assign img[14996] = 174;
assign img[14997] = 170;
assign img[14998] = 200;
assign img[14999] = 253;
assign img[15000] = 255;
assign img[15001] = 205;
assign img[15002] = 236;
assign img[15003] = 238;
assign img[15004] = 222;
assign img[15005] = 252;
assign img[15006] = 238;
assign img[15007] = 159;
assign img[15008] = 137;
assign img[15009] = 204;
assign img[15010] = 236;
assign img[15011] = 238;
assign img[15012] = 254;
assign img[15013] = 255;
assign img[15014] = 187;
assign img[15015] = 251;
assign img[15016] = 127;
assign img[15017] = 255;
assign img[15018] = 159;
assign img[15019] = 205;
assign img[15020] = 172;
assign img[15021] = 171;
assign img[15022] = 238;
assign img[15023] = 239;
assign img[15024] = 238;
assign img[15025] = 239;
assign img[15026] = 238;
assign img[15027] = 191;
assign img[15028] = 171;
assign img[15029] = 186;
assign img[15030] = 251;
assign img[15031] = 255;
assign img[15032] = 174;
assign img[15033] = 187;
assign img[15034] = 170;
assign img[15035] = 170;
assign img[15036] = 234;
assign img[15037] = 255;
assign img[15038] = 153;
assign img[15039] = 251;
assign img[15040] = 255;
assign img[15041] = 191;
assign img[15042] = 154;
assign img[15043] = 251;
assign img[15044] = 187;
assign img[15045] = 187;
assign img[15046] = 171;
assign img[15047] = 187;
assign img[15048] = 203;
assign img[15049] = 204;
assign img[15050] = 204;
assign img[15051] = 205;
assign img[15052] = 172;
assign img[15053] = 238;
assign img[15054] = 204;
assign img[15055] = 238;
assign img[15056] = 238;
assign img[15057] = 238;
assign img[15058] = 174;
assign img[15059] = 187;
assign img[15060] = 187;
assign img[15061] = 191;
assign img[15062] = 255;
assign img[15063] = 255;
assign img[15064] = 255;
assign img[15065] = 255;
assign img[15066] = 251;
assign img[15067] = 255;
assign img[15068] = 255;
assign img[15069] = 223;
assign img[15070] = 221;
assign img[15071] = 223;
assign img[15072] = 204;
assign img[15073] = 255;
assign img[15074] = 255;
assign img[15075] = 239;
assign img[15076] = 238;
assign img[15077] = 254;
assign img[15078] = 139;
assign img[15079] = 152;
assign img[15080] = 153;
assign img[15081] = 239;
assign img[15082] = 254;
assign img[15083] = 191;
assign img[15084] = 139;
assign img[15085] = 187;
assign img[15086] = 155;
assign img[15087] = 253;
assign img[15088] = 255;
assign img[15089] = 255;
assign img[15090] = 221;
assign img[15091] = 221;
assign img[15092] = 221;
assign img[15093] = 223;
assign img[15094] = 253;
assign img[15095] = 255;
assign img[15096] = 255;
assign img[15097] = 255;
assign img[15098] = 223;
assign img[15099] = 157;
assign img[15100] = 221;
assign img[15101] = 253;
assign img[15102] = 255;
assign img[15103] = 255;
assign img[15104] = 96;
assign img[15105] = 230;
assign img[15106] = 254;
assign img[15107] = 239;
assign img[15108] = 254;
assign img[15109] = 255;
assign img[15110] = 223;
assign img[15111] = 255;
assign img[15112] = 255;
assign img[15113] = 255;
assign img[15114] = 255;
assign img[15115] = 223;
assign img[15116] = 221;
assign img[15117] = 221;
assign img[15118] = 221;
assign img[15119] = 255;
assign img[15120] = 204;
assign img[15121] = 172;
assign img[15122] = 170;
assign img[15123] = 174;
assign img[15124] = 136;
assign img[15125] = 238;
assign img[15126] = 254;
assign img[15127] = 255;
assign img[15128] = 239;
assign img[15129] = 206;
assign img[15130] = 252;
assign img[15131] = 239;
assign img[15132] = 206;
assign img[15133] = 236;
assign img[15134] = 206;
assign img[15135] = 204;
assign img[15136] = 136;
assign img[15137] = 236;
assign img[15138] = 190;
assign img[15139] = 187;
assign img[15140] = 187;
assign img[15141] = 219;
assign img[15142] = 253;
assign img[15143] = 159;
assign img[15144] = 253;
assign img[15145] = 255;
assign img[15146] = 255;
assign img[15147] = 239;
assign img[15148] = 238;
assign img[15149] = 170;
assign img[15150] = 234;
assign img[15151] = 191;
assign img[15152] = 251;
assign img[15153] = 255;
assign img[15154] = 221;
assign img[15155] = 157;
assign img[15156] = 187;
assign img[15157] = 255;
assign img[15158] = 255;
assign img[15159] = 223;
assign img[15160] = 221;
assign img[15161] = 237;
assign img[15162] = 238;
assign img[15163] = 136;
assign img[15164] = 200;
assign img[15165] = 222;
assign img[15166] = 137;
assign img[15167] = 236;
assign img[15168] = 238;
assign img[15169] = 206;
assign img[15170] = 206;
assign img[15171] = 204;
assign img[15172] = 204;
assign img[15173] = 204;
assign img[15174] = 136;
assign img[15175] = 202;
assign img[15176] = 236;
assign img[15177] = 238;
assign img[15178] = 254;
assign img[15179] = 239;
assign img[15180] = 254;
assign img[15181] = 255;
assign img[15182] = 255;
assign img[15183] = 255;
assign img[15184] = 191;
assign img[15185] = 255;
assign img[15186] = 239;
assign img[15187] = 238;
assign img[15188] = 206;
assign img[15189] = 204;
assign img[15190] = 204;
assign img[15191] = 238;
assign img[15192] = 142;
assign img[15193] = 136;
assign img[15194] = 200;
assign img[15195] = 140;
assign img[15196] = 184;
assign img[15197] = 187;
assign img[15198] = 251;
assign img[15199] = 223;
assign img[15200] = 236;
assign img[15201] = 206;
assign img[15202] = 236;
assign img[15203] = 223;
assign img[15204] = 253;
assign img[15205] = 191;
assign img[15206] = 219;
assign img[15207] = 207;
assign img[15208] = 238;
assign img[15209] = 223;
assign img[15210] = 253;
assign img[15211] = 255;
assign img[15212] = 223;
assign img[15213] = 255;
assign img[15214] = 191;
assign img[15215] = 155;
assign img[15216] = 136;
assign img[15217] = 157;
assign img[15218] = 153;
assign img[15219] = 255;
assign img[15220] = 255;
assign img[15221] = 239;
assign img[15222] = 238;
assign img[15223] = 238;
assign img[15224] = 238;
assign img[15225] = 238;
assign img[15226] = 204;
assign img[15227] = 238;
assign img[15228] = 238;
assign img[15229] = 254;
assign img[15230] = 223;
assign img[15231] = 255;
assign img[15232] = 96;
assign img[15233] = 222;
assign img[15234] = 253;
assign img[15235] = 255;
assign img[15236] = 238;
assign img[15237] = 238;
assign img[15238] = 238;
assign img[15239] = 254;
assign img[15240] = 223;
assign img[15241] = 255;
assign img[15242] = 255;
assign img[15243] = 255;
assign img[15244] = 255;
assign img[15245] = 255;
assign img[15246] = 175;
assign img[15247] = 159;
assign img[15248] = 137;
assign img[15249] = 156;
assign img[15250] = 253;
assign img[15251] = 255;
assign img[15252] = 155;
assign img[15253] = 153;
assign img[15254] = 201;
assign img[15255] = 221;
assign img[15256] = 253;
assign img[15257] = 223;
assign img[15258] = 205;
assign img[15259] = 204;
assign img[15260] = 204;
assign img[15261] = 236;
assign img[15262] = 190;
assign img[15263] = 157;
assign img[15264] = 205;
assign img[15265] = 236;
assign img[15266] = 254;
assign img[15267] = 255;
assign img[15268] = 191;
assign img[15269] = 187;
assign img[15270] = 202;
assign img[15271] = 221;
assign img[15272] = 221;
assign img[15273] = 253;
assign img[15274] = 191;
assign img[15275] = 155;
assign img[15276] = 201;
assign img[15277] = 236;
assign img[15278] = 238;
assign img[15279] = 255;
assign img[15280] = 255;
assign img[15281] = 255;
assign img[15282] = 255;
assign img[15283] = 255;
assign img[15284] = 255;
assign img[15285] = 239;
assign img[15286] = 238;
assign img[15287] = 238;
assign img[15288] = 254;
assign img[15289] = 255;
assign img[15290] = 238;
assign img[15291] = 238;
assign img[15292] = 204;
assign img[15293] = 204;
assign img[15294] = 204;
assign img[15295] = 204;
assign img[15296] = 220;
assign img[15297] = 221;
assign img[15298] = 221;
assign img[15299] = 253;
assign img[15300] = 223;
assign img[15301] = 221;
assign img[15302] = 137;
assign img[15303] = 136;
assign img[15304] = 184;
assign img[15305] = 155;
assign img[15306] = 217;
assign img[15307] = 239;
assign img[15308] = 238;
assign img[15309] = 238;
assign img[15310] = 220;
assign img[15311] = 221;
assign img[15312] = 253;
assign img[15313] = 255;
assign img[15314] = 255;
assign img[15315] = 223;
assign img[15316] = 221;
assign img[15317] = 221;
assign img[15318] = 253;
assign img[15319] = 223;
assign img[15320] = 221;
assign img[15321] = 221;
assign img[15322] = 237;
assign img[15323] = 238;
assign img[15324] = 238;
assign img[15325] = 238;
assign img[15326] = 238;
assign img[15327] = 223;
assign img[15328] = 204;
assign img[15329] = 204;
assign img[15330] = 236;
assign img[15331] = 223;
assign img[15332] = 221;
assign img[15333] = 221;
assign img[15334] = 157;
assign img[15335] = 185;
assign img[15336] = 187;
assign img[15337] = 255;
assign img[15338] = 255;
assign img[15339] = 255;
assign img[15340] = 140;
assign img[15341] = 238;
assign img[15342] = 238;
assign img[15343] = 223;
assign img[15344] = 204;
assign img[15345] = 238;
assign img[15346] = 187;
assign img[15347] = 239;
assign img[15348] = 254;
assign img[15349] = 255;
assign img[15350] = 255;
assign img[15351] = 255;
assign img[15352] = 255;
assign img[15353] = 239;
assign img[15354] = 238;
assign img[15355] = 207;
assign img[15356] = 204;
assign img[15357] = 253;
assign img[15358] = 223;
assign img[15359] = 253;
assign img[15360] = 96;
assign img[15361] = 206;
assign img[15362] = 236;
assign img[15363] = 238;
assign img[15364] = 238;
assign img[15365] = 238;
assign img[15366] = 254;
assign img[15367] = 255;
assign img[15368] = 239;
assign img[15369] = 238;
assign img[15370] = 238;
assign img[15371] = 174;
assign img[15372] = 170;
assign img[15373] = 238;
assign img[15374] = 206;
assign img[15375] = 204;
assign img[15376] = 236;
assign img[15377] = 206;
assign img[15378] = 236;
assign img[15379] = 255;
assign img[15380] = 170;
assign img[15381] = 238;
assign img[15382] = 174;
assign img[15383] = 238;
assign img[15384] = 238;
assign img[15385] = 255;
assign img[15386] = 171;
assign img[15387] = 251;
assign img[15388] = 251;
assign img[15389] = 255;
assign img[15390] = 223;
assign img[15391] = 205;
assign img[15392] = 185;
assign img[15393] = 187;
assign img[15394] = 171;
assign img[15395] = 170;
assign img[15396] = 187;
assign img[15397] = 255;
assign img[15398] = 255;
assign img[15399] = 255;
assign img[15400] = 221;
assign img[15401] = 221;
assign img[15402] = 238;
assign img[15403] = 255;
assign img[15404] = 187;
assign img[15405] = 171;
assign img[15406] = 238;
assign img[15407] = 174;
assign img[15408] = 234;
assign img[15409] = 255;
assign img[15410] = 255;
assign img[15411] = 191;
assign img[15412] = 187;
assign img[15413] = 255;
assign img[15414] = 223;
assign img[15415] = 223;
assign img[15416] = 253;
assign img[15417] = 205;
assign img[15418] = 172;
assign img[15419] = 170;
assign img[15420] = 234;
assign img[15421] = 191;
assign img[15422] = 251;
assign img[15423] = 255;
assign img[15424] = 238;
assign img[15425] = 206;
assign img[15426] = 236;
assign img[15427] = 238;
assign img[15428] = 206;
assign img[15429] = 157;
assign img[15430] = 137;
assign img[15431] = 136;
assign img[15432] = 200;
assign img[15433] = 204;
assign img[15434] = 236;
assign img[15435] = 238;
assign img[15436] = 238;
assign img[15437] = 238;
assign img[15438] = 238;
assign img[15439] = 238;
assign img[15440] = 190;
assign img[15441] = 254;
assign img[15442] = 255;
assign img[15443] = 238;
assign img[15444] = 204;
assign img[15445] = 221;
assign img[15446] = 137;
assign img[15447] = 236;
assign img[15448] = 254;
assign img[15449] = 221;
assign img[15450] = 205;
assign img[15451] = 252;
assign img[15452] = 206;
assign img[15453] = 204;
assign img[15454] = 252;
assign img[15455] = 191;
assign img[15456] = 187;
assign img[15457] = 155;
assign img[15458] = 250;
assign img[15459] = 255;
assign img[15460] = 238;
assign img[15461] = 170;
assign img[15462] = 170;
assign img[15463] = 251;
assign img[15464] = 255;
assign img[15465] = 255;
assign img[15466] = 255;
assign img[15467] = 255;
assign img[15468] = 238;
assign img[15469] = 238;
assign img[15470] = 222;
assign img[15471] = 255;
assign img[15472] = 223;
assign img[15473] = 221;
assign img[15474] = 236;
assign img[15475] = 255;
assign img[15476] = 191;
assign img[15477] = 187;
assign img[15478] = 234;
assign img[15479] = 255;
assign img[15480] = 238;
assign img[15481] = 255;
assign img[15482] = 255;
assign img[15483] = 255;
assign img[15484] = 255;
assign img[15485] = 255;
assign img[15486] = 223;
assign img[15487] = 255;
assign img[15488] = 96;
assign img[15489] = 206;
assign img[15490] = 252;
assign img[15491] = 175;
assign img[15492] = 170;
assign img[15493] = 238;
assign img[15494] = 238;
assign img[15495] = 191;
assign img[15496] = 251;
assign img[15497] = 255;
assign img[15498] = 255;
assign img[15499] = 255;
assign img[15500] = 238;
assign img[15501] = 254;
assign img[15502] = 223;
assign img[15503] = 221;
assign img[15504] = 204;
assign img[15505] = 221;
assign img[15506] = 236;
assign img[15507] = 238;
assign img[15508] = 238;
assign img[15509] = 238;
assign img[15510] = 238;
assign img[15511] = 255;
assign img[15512] = 255;
assign img[15513] = 255;
assign img[15514] = 255;
assign img[15515] = 255;
assign img[15516] = 238;
assign img[15517] = 238;
assign img[15518] = 238;
assign img[15519] = 238;
assign img[15520] = 170;
assign img[15521] = 234;
assign img[15522] = 238;
assign img[15523] = 238;
assign img[15524] = 238;
assign img[15525] = 206;
assign img[15526] = 221;
assign img[15527] = 157;
assign img[15528] = 217;
assign img[15529] = 205;
assign img[15530] = 236;
assign img[15531] = 254;
assign img[15532] = 223;
assign img[15533] = 205;
assign img[15534] = 236;
assign img[15535] = 255;
assign img[15536] = 255;
assign img[15537] = 255;
assign img[15538] = 255;
assign img[15539] = 255;
assign img[15540] = 255;
assign img[15541] = 255;
assign img[15542] = 255;
assign img[15543] = 255;
assign img[15544] = 223;
assign img[15545] = 205;
assign img[15546] = 140;
assign img[15547] = 186;
assign img[15548] = 255;
assign img[15549] = 255;
assign img[15550] = 255;
assign img[15551] = 255;
assign img[15552] = 238;
assign img[15553] = 254;
assign img[15554] = 255;
assign img[15555] = 255;
assign img[15556] = 207;
assign img[15557] = 255;
assign img[15558] = 155;
assign img[15559] = 221;
assign img[15560] = 221;
assign img[15561] = 223;
assign img[15562] = 221;
assign img[15563] = 221;
assign img[15564] = 221;
assign img[15565] = 223;
assign img[15566] = 205;
assign img[15567] = 238;
assign img[15568] = 238;
assign img[15569] = 238;
assign img[15570] = 238;
assign img[15571] = 238;
assign img[15572] = 204;
assign img[15573] = 236;
assign img[15574] = 170;
assign img[15575] = 186;
assign img[15576] = 217;
assign img[15577] = 191;
assign img[15578] = 238;
assign img[15579] = 255;
assign img[15580] = 238;
assign img[15581] = 238;
assign img[15582] = 238;
assign img[15583] = 175;
assign img[15584] = 234;
assign img[15585] = 138;
assign img[15586] = 238;
assign img[15587] = 239;
assign img[15588] = 238;
assign img[15589] = 254;
assign img[15590] = 255;
assign img[15591] = 255;
assign img[15592] = 255;
assign img[15593] = 255;
assign img[15594] = 255;
assign img[15595] = 255;
assign img[15596] = 255;
assign img[15597] = 255;
assign img[15598] = 223;
assign img[15599] = 223;
assign img[15600] = 207;
assign img[15601] = 206;
assign img[15602] = 238;
assign img[15603] = 255;
assign img[15604] = 238;
assign img[15605] = 238;
assign img[15606] = 238;
assign img[15607] = 238;
assign img[15608] = 238;
assign img[15609] = 255;
assign img[15610] = 255;
assign img[15611] = 239;
assign img[15612] = 238;
assign img[15613] = 254;
assign img[15614] = 255;
assign img[15615] = 255;
assign img[15616] = 64;
assign img[15617] = 204;
assign img[15618] = 236;
assign img[15619] = 238;
assign img[15620] = 238;
assign img[15621] = 238;
assign img[15622] = 222;
assign img[15623] = 255;
assign img[15624] = 255;
assign img[15625] = 255;
assign img[15626] = 220;
assign img[15627] = 255;
assign img[15628] = 255;
assign img[15629] = 255;
assign img[15630] = 255;
assign img[15631] = 223;
assign img[15632] = 205;
assign img[15633] = 204;
assign img[15634] = 236;
assign img[15635] = 174;
assign img[15636] = 138;
assign img[15637] = 255;
assign img[15638] = 255;
assign img[15639] = 239;
assign img[15640] = 238;
assign img[15641] = 238;
assign img[15642] = 254;
assign img[15643] = 255;
assign img[15644] = 255;
assign img[15645] = 255;
assign img[15646] = 238;
assign img[15647] = 255;
assign img[15648] = 63;
assign img[15649] = 247;
assign img[15650] = 223;
assign img[15651] = 255;
assign img[15652] = 255;
assign img[15653] = 191;
assign img[15654] = 187;
assign img[15655] = 187;
assign img[15656] = 234;
assign img[15657] = 254;
assign img[15658] = 255;
assign img[15659] = 255;
assign img[15660] = 251;
assign img[15661] = 255;
assign img[15662] = 238;
assign img[15663] = 191;
assign img[15664] = 187;
assign img[15665] = 255;
assign img[15666] = 255;
assign img[15667] = 255;
assign img[15668] = 157;
assign img[15669] = 255;
assign img[15670] = 255;
assign img[15671] = 255;
assign img[15672] = 255;
assign img[15673] = 255;
assign img[15674] = 255;
assign img[15675] = 255;
assign img[15676] = 187;
assign img[15677] = 239;
assign img[15678] = 238;
assign img[15679] = 254;
assign img[15680] = 255;
assign img[15681] = 255;
assign img[15682] = 221;
assign img[15683] = 237;
assign img[15684] = 238;
assign img[15685] = 206;
assign img[15686] = 220;
assign img[15687] = 253;
assign img[15688] = 159;
assign img[15689] = 153;
assign img[15690] = 232;
assign img[15691] = 174;
assign img[15692] = 234;
assign img[15693] = 238;
assign img[15694] = 238;
assign img[15695] = 254;
assign img[15696] = 255;
assign img[15697] = 255;
assign img[15698] = 239;
assign img[15699] = 238;
assign img[15700] = 170;
assign img[15701] = 170;
assign img[15702] = 234;
assign img[15703] = 238;
assign img[15704] = 174;
assign img[15705] = 186;
assign img[15706] = 170;
assign img[15707] = 170;
assign img[15708] = 234;
assign img[15709] = 238;
assign img[15710] = 238;
assign img[15711] = 174;
assign img[15712] = 234;
assign img[15713] = 191;
assign img[15714] = 171;
assign img[15715] = 190;
assign img[15716] = 187;
assign img[15717] = 255;
assign img[15718] = 238;
assign img[15719] = 238;
assign img[15720] = 238;
assign img[15721] = 254;
assign img[15722] = 255;
assign img[15723] = 223;
assign img[15724] = 153;
assign img[15725] = 255;
assign img[15726] = 255;
assign img[15727] = 255;
assign img[15728] = 255;
assign img[15729] = 255;
assign img[15730] = 255;
assign img[15731] = 255;
assign img[15732] = 255;
assign img[15733] = 255;
assign img[15734] = 223;
assign img[15735] = 255;
assign img[15736] = 255;
assign img[15737] = 255;
assign img[15738] = 255;
assign img[15739] = 255;
assign img[15740] = 255;
assign img[15741] = 255;
assign img[15742] = 255;
assign img[15743] = 223;
assign img[15744] = 96;
assign img[15745] = 238;
assign img[15746] = 254;
assign img[15747] = 255;
assign img[15748] = 238;
assign img[15749] = 238;
assign img[15750] = 206;
assign img[15751] = 204;
assign img[15752] = 236;
assign img[15753] = 238;
assign img[15754] = 238;
assign img[15755] = 174;
assign img[15756] = 238;
assign img[15757] = 255;
assign img[15758] = 255;
assign img[15759] = 223;
assign img[15760] = 253;
assign img[15761] = 255;
assign img[15762] = 238;
assign img[15763] = 255;
assign img[15764] = 238;
assign img[15765] = 238;
assign img[15766] = 238;
assign img[15767] = 255;
assign img[15768] = 238;
assign img[15769] = 255;
assign img[15770] = 127;
assign img[15771] = 239;
assign img[15772] = 206;
assign img[15773] = 238;
assign img[15774] = 206;
assign img[15775] = 156;
assign img[15776] = 185;
assign img[15777] = 251;
assign img[15778] = 223;
assign img[15779] = 255;
assign img[15780] = 239;
assign img[15781] = 238;
assign img[15782] = 206;
assign img[15783] = 207;
assign img[15784] = 238;
assign img[15785] = 223;
assign img[15786] = 157;
assign img[15787] = 153;
assign img[15788] = 201;
assign img[15789] = 204;
assign img[15790] = 236;
assign img[15791] = 238;
assign img[15792] = 204;
assign img[15793] = 220;
assign img[15794] = 221;
assign img[15795] = 255;
assign img[15796] = 255;
assign img[15797] = 223;
assign img[15798] = 221;
assign img[15799] = 223;
assign img[15800] = 255;
assign img[15801] = 205;
assign img[15802] = 204;
assign img[15803] = 205;
assign img[15804] = 236;
assign img[15805] = 255;
assign img[15806] = 187;
assign img[15807] = 255;
assign img[15808] = 255;
assign img[15809] = 239;
assign img[15810] = 238;
assign img[15811] = 238;
assign img[15812] = 206;
assign img[15813] = 190;
assign img[15814] = 255;
assign img[15815] = 239;
assign img[15816] = 206;
assign img[15817] = 204;
assign img[15818] = 204;
assign img[15819] = 189;
assign img[15820] = 251;
assign img[15821] = 143;
assign img[15822] = 204;
assign img[15823] = 236;
assign img[15824] = 238;
assign img[15825] = 238;
assign img[15826] = 238;
assign img[15827] = 238;
assign img[15828] = 174;
assign img[15829] = 170;
assign img[15830] = 234;
assign img[15831] = 238;
assign img[15832] = 206;
assign img[15833] = 221;
assign img[15834] = 205;
assign img[15835] = 204;
assign img[15836] = 236;
assign img[15837] = 206;
assign img[15838] = 236;
assign img[15839] = 191;
assign img[15840] = 187;
assign img[15841] = 219;
assign img[15842] = 236;
assign img[15843] = 255;
assign img[15844] = 221;
assign img[15845] = 239;
assign img[15846] = 238;
assign img[15847] = 238;
assign img[15848] = 238;
assign img[15849] = 254;
assign img[15850] = 187;
assign img[15851] = 255;
assign img[15852] = 255;
assign img[15853] = 255;
assign img[15854] = 255;
assign img[15855] = 239;
assign img[15856] = 254;
assign img[15857] = 239;
assign img[15858] = 254;
assign img[15859] = 255;
assign img[15860] = 191;
assign img[15861] = 171;
assign img[15862] = 234;
assign img[15863] = 238;
assign img[15864] = 254;
assign img[15865] = 223;
assign img[15866] = 221;
assign img[15867] = 221;
assign img[15868] = 236;
assign img[15869] = 254;
assign img[15870] = 239;
assign img[15871] = 255;
assign img[15872] = 64;
assign img[15873] = 213;
assign img[15874] = 253;
assign img[15875] = 223;
assign img[15876] = 141;
assign img[15877] = 238;
assign img[15878] = 238;
assign img[15879] = 238;
assign img[15880] = 238;
assign img[15881] = 238;
assign img[15882] = 222;
assign img[15883] = 223;
assign img[15884] = 221;
assign img[15885] = 221;
assign img[15886] = 221;
assign img[15887] = 221;
assign img[15888] = 221;
assign img[15889] = 253;
assign img[15890] = 255;
assign img[15891] = 255;
assign img[15892] = 255;
assign img[15893] = 255;
assign img[15894] = 255;
assign img[15895] = 255;
assign img[15896] = 255;
assign img[15897] = 191;
assign img[15898] = 187;
assign img[15899] = 187;
assign img[15900] = 187;
assign img[15901] = 187;
assign img[15902] = 255;
assign img[15903] = 191;
assign img[15904] = 170;
assign img[15905] = 170;
assign img[15906] = 202;
assign img[15907] = 238;
assign img[15908] = 222;
assign img[15909] = 221;
assign img[15910] = 205;
assign img[15911] = 220;
assign img[15912] = 221;
assign img[15913] = 221;
assign img[15914] = 221;
assign img[15915] = 205;
assign img[15916] = 220;
assign img[15917] = 141;
assign img[15918] = 153;
assign img[15919] = 171;
assign img[15920] = 250;
assign img[15921] = 255;
assign img[15922] = 255;
assign img[15923] = 223;
assign img[15924] = 189;
assign img[15925] = 255;
assign img[15926] = 255;
assign img[15927] = 239;
assign img[15928] = 174;
assign img[15929] = 170;
assign img[15930] = 234;
assign img[15931] = 238;
assign img[15932] = 254;
assign img[15933] = 191;
assign img[15934] = 223;
assign img[15935] = 255;
assign img[15936] = 255;
assign img[15937] = 255;
assign img[15938] = 221;
assign img[15939] = 255;
assign img[15940] = 239;
assign img[15941] = 238;
assign img[15942] = 220;
assign img[15943] = 157;
assign img[15944] = 249;
assign img[15945] = 255;
assign img[15946] = 238;
assign img[15947] = 191;
assign img[15948] = 170;
assign img[15949] = 154;
assign img[15950] = 249;
assign img[15951] = 255;
assign img[15952] = 255;
assign img[15953] = 255;
assign img[15954] = 175;
assign img[15955] = 238;
assign img[15956] = 206;
assign img[15957] = 238;
assign img[15958] = 206;
assign img[15959] = 204;
assign img[15960] = 204;
assign img[15961] = 221;
assign img[15962] = 204;
assign img[15963] = 204;
assign img[15964] = 236;
assign img[15965] = 238;
assign img[15966] = 254;
assign img[15967] = 255;
assign img[15968] = 171;
assign img[15969] = 170;
assign img[15970] = 234;
assign img[15971] = 238;
assign img[15972] = 238;
assign img[15973] = 238;
assign img[15974] = 238;
assign img[15975] = 238;
assign img[15976] = 254;
assign img[15977] = 255;
assign img[15978] = 255;
assign img[15979] = 239;
assign img[15980] = 206;
assign img[15981] = 238;
assign img[15982] = 254;
assign img[15983] = 223;
assign img[15984] = 221;
assign img[15985] = 221;
assign img[15986] = 221;
assign img[15987] = 221;
assign img[15988] = 221;
assign img[15989] = 221;
assign img[15990] = 253;
assign img[15991] = 255;
assign img[15992] = 255;
assign img[15993] = 255;
assign img[15994] = 238;
assign img[15995] = 255;
assign img[15996] = 238;
assign img[15997] = 255;
assign img[15998] = 255;
assign img[15999] = 255;
assign img[16000] = 112;
assign img[16001] = 255;
assign img[16002] = 255;
assign img[16003] = 255;
assign img[16004] = 205;
assign img[16005] = 221;
assign img[16006] = 221;
assign img[16007] = 253;
assign img[16008] = 255;
assign img[16009] = 255;
assign img[16010] = 223;
assign img[16011] = 221;
assign img[16012] = 221;
assign img[16013] = 253;
assign img[16014] = 159;
assign img[16015] = 187;
assign img[16016] = 187;
assign img[16017] = 187;
assign img[16018] = 251;
assign img[16019] = 255;
assign img[16020] = 204;
assign img[16021] = 236;
assign img[16022] = 206;
assign img[16023] = 236;
assign img[16024] = 238;
assign img[16025] = 239;
assign img[16026] = 238;
assign img[16027] = 255;
assign img[16028] = 223;
assign img[16029] = 255;
assign img[16030] = 239;
assign img[16031] = 238;
assign img[16032] = 138;
assign img[16033] = 238;
assign img[16034] = 206;
assign img[16035] = 238;
assign img[16036] = 206;
assign img[16037] = 253;
assign img[16038] = 255;
assign img[16039] = 255;
assign img[16040] = 187;
assign img[16041] = 187;
assign img[16042] = 187;
assign img[16043] = 187;
assign img[16044] = 139;
assign img[16045] = 136;
assign img[16046] = 232;
assign img[16047] = 238;
assign img[16048] = 238;
assign img[16049] = 255;
assign img[16050] = 255;
assign img[16051] = 255;
assign img[16052] = 238;
assign img[16053] = 238;
assign img[16054] = 222;
assign img[16055] = 221;
assign img[16056] = 255;
assign img[16057] = 191;
assign img[16058] = 187;
assign img[16059] = 187;
assign img[16060] = 255;
assign img[16061] = 191;
assign img[16062] = 187;
assign img[16063] = 187;
assign img[16064] = 170;
assign img[16065] = 238;
assign img[16066] = 190;
assign img[16067] = 255;
assign img[16068] = 175;
assign img[16069] = 170;
assign img[16070] = 170;
assign img[16071] = 170;
assign img[16072] = 202;
assign img[16073] = 204;
assign img[16074] = 236;
assign img[16075] = 238;
assign img[16076] = 170;
assign img[16077] = 255;
assign img[16078] = 204;
assign img[16079] = 253;
assign img[16080] = 255;
assign img[16081] = 255;
assign img[16082] = 254;
assign img[16083] = 223;
assign img[16084] = 172;
assign img[16085] = 170;
assign img[16086] = 170;
assign img[16087] = 170;
assign img[16088] = 170;
assign img[16089] = 170;
assign img[16090] = 238;
assign img[16091] = 206;
assign img[16092] = 238;
assign img[16093] = 206;
assign img[16094] = 236;
assign img[16095] = 207;
assign img[16096] = 236;
assign img[16097] = 238;
assign img[16098] = 238;
assign img[16099] = 255;
assign img[16100] = 221;
assign img[16101] = 255;
assign img[16102] = 205;
assign img[16103] = 236;
assign img[16104] = 238;
assign img[16105] = 220;
assign img[16106] = 253;
assign img[16107] = 223;
assign img[16108] = 204;
assign img[16109] = 220;
assign img[16110] = 221;
assign img[16111] = 221;
assign img[16112] = 221;
assign img[16113] = 157;
assign img[16114] = 185;
assign img[16115] = 223;
assign img[16116] = 221;
assign img[16117] = 205;
assign img[16118] = 236;
assign img[16119] = 238;
assign img[16120] = 238;
assign img[16121] = 238;
assign img[16122] = 220;
assign img[16123] = 205;
assign img[16124] = 204;
assign img[16125] = 236;
assign img[16126] = 238;
assign img[16127] = 238;
assign img[16128] = 0;
assign img[16129] = 145;
assign img[16130] = 249;
assign img[16131] = 255;
assign img[16132] = 206;
assign img[16133] = 236;
assign img[16134] = 206;
assign img[16135] = 252;
assign img[16136] = 238;
assign img[16137] = 255;
assign img[16138] = 255;
assign img[16139] = 255;
assign img[16140] = 255;
assign img[16141] = 255;
assign img[16142] = 255;
assign img[16143] = 239;
assign img[16144] = 238;
assign img[16145] = 254;
assign img[16146] = 239;
assign img[16147] = 206;
assign img[16148] = 236;
assign img[16149] = 238;
assign img[16150] = 238;
assign img[16151] = 238;
assign img[16152] = 255;
assign img[16153] = 239;
assign img[16154] = 254;
assign img[16155] = 223;
assign img[16156] = 255;
assign img[16157] = 255;
assign img[16158] = 207;
assign img[16159] = 205;
assign img[16160] = 136;
assign img[16161] = 170;
assign img[16162] = 138;
assign img[16163] = 136;
assign img[16164] = 136;
assign img[16165] = 236;
assign img[16166] = 238;
assign img[16167] = 238;
assign img[16168] = 238;
assign img[16169] = 222;
assign img[16170] = 221;
assign img[16171] = 207;
assign img[16172] = 204;
assign img[16173] = 204;
assign img[16174] = 236;
assign img[16175] = 238;
assign img[16176] = 238;
assign img[16177] = 206;
assign img[16178] = 204;
assign img[16179] = 204;
assign img[16180] = 204;
assign img[16181] = 252;
assign img[16182] = 206;
assign img[16183] = 238;
assign img[16184] = 204;
assign img[16185] = 238;
assign img[16186] = 204;
assign img[16187] = 206;
assign img[16188] = 254;
assign img[16189] = 159;
assign img[16190] = 221;
assign img[16191] = 252;
assign img[16192] = 238;
assign img[16193] = 238;
assign img[16194] = 220;
assign img[16195] = 253;
assign img[16196] = 223;
assign img[16197] = 221;
assign img[16198] = 221;
assign img[16199] = 221;
assign img[16200] = 221;
assign img[16201] = 255;
assign img[16202] = 238;
assign img[16203] = 238;
assign img[16204] = 206;
assign img[16205] = 206;
assign img[16206] = 252;
assign img[16207] = 255;
assign img[16208] = 255;
assign img[16209] = 255;
assign img[16210] = 255;
assign img[16211] = 255;
assign img[16212] = 255;
assign img[16213] = 255;
assign img[16214] = 154;
assign img[16215] = 223;
assign img[16216] = 205;
assign img[16217] = 238;
assign img[16218] = 238;
assign img[16219] = 255;
assign img[16220] = 236;
assign img[16221] = 238;
assign img[16222] = 238;
assign img[16223] = 174;
assign img[16224] = 170;
assign img[16225] = 238;
assign img[16226] = 238;
assign img[16227] = 238;
assign img[16228] = 220;
assign img[16229] = 221;
assign img[16230] = 153;
assign img[16231] = 217;
assign img[16232] = 253;
assign img[16233] = 255;
assign img[16234] = 255;
assign img[16235] = 255;
assign img[16236] = 237;
assign img[16237] = 255;
assign img[16238] = 255;
assign img[16239] = 223;
assign img[16240] = 204;
assign img[16241] = 204;
assign img[16242] = 236;
assign img[16243] = 238;
assign img[16244] = 222;
assign img[16245] = 205;
assign img[16246] = 236;
assign img[16247] = 238;
assign img[16248] = 238;
assign img[16249] = 238;
assign img[16250] = 238;
assign img[16251] = 238;
assign img[16252] = 238;
assign img[16253] = 238;
assign img[16254] = 206;
assign img[16255] = 221;
assign img[16256] = 96;
assign img[16257] = 238;
assign img[16258] = 238;
assign img[16259] = 239;
assign img[16260] = 238;
assign img[16261] = 254;
assign img[16262] = 191;
assign img[16263] = 170;
assign img[16264] = 234;
assign img[16265] = 238;
assign img[16266] = 238;
assign img[16267] = 238;
assign img[16268] = 138;
assign img[16269] = 136;
assign img[16270] = 236;
assign img[16271] = 206;
assign img[16272] = 204;
assign img[16273] = 204;
assign img[16274] = 254;
assign img[16275] = 255;
assign img[16276] = 223;
assign img[16277] = 253;
assign img[16278] = 255;
assign img[16279] = 255;
assign img[16280] = 255;
assign img[16281] = 223;
assign img[16282] = 205;
assign img[16283] = 238;
assign img[16284] = 206;
assign img[16285] = 204;
assign img[16286] = 204;
assign img[16287] = 204;
assign img[16288] = 204;
assign img[16289] = 236;
assign img[16290] = 254;
assign img[16291] = 239;
assign img[16292] = 238;
assign img[16293] = 238;
assign img[16294] = 252;
assign img[16295] = 221;
assign img[16296] = 253;
assign img[16297] = 255;
assign img[16298] = 255;
assign img[16299] = 239;
assign img[16300] = 140;
assign img[16301] = 136;
assign img[16302] = 232;
assign img[16303] = 206;
assign img[16304] = 236;
assign img[16305] = 255;
assign img[16306] = 238;
assign img[16307] = 223;
assign img[16308] = 253;
assign img[16309] = 255;
assign img[16310] = 205;
assign img[16311] = 221;
assign img[16312] = 221;
assign img[16313] = 253;
assign img[16314] = 221;
assign img[16315] = 221;
assign img[16316] = 200;
assign img[16317] = 221;
assign img[16318] = 253;
assign img[16319] = 255;
assign img[16320] = 255;
assign img[16321] = 255;
assign img[16322] = 255;
assign img[16323] = 255;
assign img[16324] = 207;
assign img[16325] = 191;
assign img[16326] = 187;
assign img[16327] = 139;
assign img[16328] = 136;
assign img[16329] = 136;
assign img[16330] = 200;
assign img[16331] = 253;
assign img[16332] = 223;
assign img[16333] = 221;
assign img[16334] = 205;
assign img[16335] = 238;
assign img[16336] = 222;
assign img[16337] = 253;
assign img[16338] = 255;
assign img[16339] = 239;
assign img[16340] = 206;
assign img[16341] = 172;
assign img[16342] = 186;
assign img[16343] = 255;
assign img[16344] = 223;
assign img[16345] = 221;
assign img[16346] = 253;
assign img[16347] = 255;
assign img[16348] = 255;
assign img[16349] = 255;
assign img[16350] = 137;
assign img[16351] = 136;
assign img[16352] = 152;
assign img[16353] = 217;
assign img[16354] = 253;
assign img[16355] = 239;
assign img[16356] = 238;
assign img[16357] = 239;
assign img[16358] = 255;
assign img[16359] = 255;
assign img[16360] = 255;
assign img[16361] = 255;
assign img[16362] = 238;
assign img[16363] = 255;
assign img[16364] = 221;
assign img[16365] = 255;
assign img[16366] = 255;
assign img[16367] = 255;
assign img[16368] = 255;
assign img[16369] = 255;
assign img[16370] = 255;
assign img[16371] = 223;
assign img[16372] = 253;
assign img[16373] = 239;
assign img[16374] = 238;
assign img[16375] = 238;
assign img[16376] = 238;
assign img[16377] = 238;
assign img[16378] = 170;
assign img[16379] = 171;
assign img[16380] = 234;
assign img[16381] = 255;
assign img[16382] = 223;
assign img[16383] = 238;
    
endmodule
